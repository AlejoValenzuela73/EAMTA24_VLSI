magic
tech sky130A
magscale 1 2
timestamp 1709751578
<< nwell >>
rect -109 -177 109 177
<< pmos >>
rect -15 -115 15 115
<< pdiff >>
rect -73 103 -15 115
rect -73 -103 -61 103
rect -27 -103 -15 103
rect -73 -115 -15 -103
rect 15 103 73 115
rect 15 -103 27 103
rect 61 -103 73 103
rect 15 -115 73 -103
<< pdiffc >>
rect -61 -103 -27 103
rect 27 -103 61 103
<< poly >>
rect -15 115 15 141
rect -15 -141 15 -115
<< locali >>
rect -61 103 -27 119
rect -61 -119 -27 -103
rect 27 103 61 119
rect 27 -119 61 -103
<< viali >>
rect -61 -103 -27 103
rect 27 -103 61 103
<< metal1 >>
rect -67 103 -21 115
rect -67 -103 -61 103
rect -27 -103 -21 103
rect -67 -115 -21 -103
rect 21 103 67 115
rect 21 -103 27 103
rect 61 -103 67 103
rect 21 -115 67 -103
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.15 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
