magic
tech sky130A
timestamp 1710544241
use bctr  bctr_0 bitcounter
timestamp 1710544241
transform 1 0 852 0 1 3
box -852 -3 1473 541
<< end >>
