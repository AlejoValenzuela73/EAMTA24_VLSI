magic
tech sky130A
magscale 1 2
timestamp 1709826131
use grid  grid_0
timestamp 1678218586
transform 1 0 61 0 1 10
box -61 -10 259 1053
use sky130_fd_pr__nfet_01v8_5CZXLZ  sky130_fd_pr__nfet_01v8_5CZXLZ_0
timestamp 1709826131
transform 1 0 526 0 1 664
box -73 -101 73 101
use sky130_fd_pr__nfet_01v8_5CZXLZ  sky130_fd_pr__nfet_01v8_5CZXLZ_1
timestamp 1709826131
transform 1 0 -155 0 1 217
box -73 -101 73 101
use sky130_fd_pr__pfet_01v8_5EUKDE  sky130_fd_pr__pfet_01v8_5EUKDE_0
timestamp 1709826131
transform 1 0 246 0 1 627
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_5EUKDE  sky130_fd_pr__pfet_01v8_5EUKDE_1
timestamp 1709826131
transform 1 0 158 0 1 627
box -109 -362 109 362
<< end >>
