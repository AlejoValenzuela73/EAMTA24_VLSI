magic
tech sky130A
magscale 1 2
timestamp 1710535082
<< nwell >>
rect -78 1074 290 1082
rect -78 1070 306 1074
rect -78 1068 304 1070
rect -1054 1034 -933 1064
rect -1054 1016 -640 1034
rect -1054 990 -784 1016
rect -1054 972 -933 990
rect -1054 964 -942 972
rect -1054 886 -916 964
rect -868 886 -860 964
rect -1054 876 -940 886
rect -1054 511 -933 876
rect -14 556 304 1068
rect -16 520 994 556
rect -16 519 274 520
rect -20 514 274 519
rect -1054 494 -888 511
rect -975 484 -888 494
rect -22 508 274 514
rect 420 508 994 520
rect -22 496 218 508
rect -22 490 280 496
rect 512 490 994 508
rect 512 482 698 490
<< metal1 >>
rect -1008 1024 -640 1034
rect -1030 1016 -640 1024
rect -1030 994 -946 1016
rect -934 954 -860 964
rect -934 892 -930 954
rect -866 892 -860 954
rect -934 886 -860 892
rect -1014 4 -621 52
rect -47 4 135 55
<< via1 >>
rect -930 892 -866 954
<< metal2 >>
rect -950 954 -846 966
rect -950 892 -930 954
rect -866 892 -846 954
rect -950 878 -846 892
rect 0 508 70 624
rect -104 436 72 508
rect 12 310 50 312
rect 10 294 50 310
rect -1666 292 50 294
rect -1666 244 52 292
rect -1656 230 52 244
rect -1656 220 50 230
rect -1656 218 18 220
use and  and_0 and
timestamp 1709929695
transform 1 0 -1607 0 1 -1
box -6 0 632 1063
use ffdr3  ffdr3_0 ffdr
timestamp 1710534732
transform 1 0 322 0 1 2
box -322 -2 2624 1079
use xor  xor_0 xor
timestamp 1710533398
transform 1 0 -662 0 1 0
box -310 -2 652 1074
<< end >>
