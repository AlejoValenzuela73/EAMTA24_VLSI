magic
tech sky130A
timestamp 1710559709
<< nwell >>
rect 8 -424 77 -414
rect 7 -449 78 -424
rect 8 -466 77 -449
rect 2222 -466 2304 -391
rect -5 -585 2304 -466
rect -5 -766 2296 -585
<< metal1 >>
rect 2 129 85 144
rect 2 88 20 129
rect 65 88 85 129
rect 2 64 85 88
rect 20 26 191 29
rect 1 -42 2322 26
rect 21 -428 92 -406
rect 21 -461 33 -428
rect 71 -461 92 -428
rect 21 -487 92 -461
rect 19 -607 2299 -518
rect 19 -609 1943 -607
rect 2098 -609 2299 -607
rect 8 -961 82 -934
rect 8 -1010 20 -961
rect 66 -1010 82 -961
rect 8 -1029 82 -1010
rect -7 -1088 299 -1072
rect 372 -1088 509 -1073
rect -7 -1090 305 -1088
rect 306 -1090 509 -1088
rect -7 -1098 509 -1090
rect 513 -1098 2311 -1082
rect -7 -1142 2311 -1098
rect -7 -1154 326 -1142
rect 331 -1149 2311 -1142
rect 11 -1157 326 -1154
<< via1 >>
rect 20 88 65 129
rect 33 -461 71 -428
rect 20 -1010 66 -961
<< metal2 >>
rect 1861 504 1919 517
rect 1861 469 1874 504
rect 1906 469 1919 504
rect 1861 459 1919 469
rect 6 129 77 132
rect 6 88 20 129
rect 65 88 77 129
rect 6 83 77 88
rect 22 -428 83 -420
rect 22 -461 33 -428
rect 71 -461 83 -428
rect 22 -469 83 -461
rect -1 -799 61 -794
rect -1 -816 66 -799
rect -1 -853 18 -816
rect 51 -853 66 -816
rect -1 -870 66 -853
rect 8 -961 82 -948
rect 8 -1010 20 -961
rect 66 -1010 82 -961
rect 8 -1024 82 -1010
rect 3 -1367 72 -1347
rect 3 -1407 18 -1367
rect 53 -1407 72 -1367
rect 3 -1410 72 -1407
<< via2 >>
rect 1874 469 1906 504
rect 20 88 65 129
rect 1493 126 1522 155
rect 1492 -167 1521 -138
rect 24 -302 54 -274
rect 34 -459 69 -430
rect 18 -853 51 -816
rect 20 -1010 66 -961
rect 18 -1407 53 -1367
<< metal3 >>
rect 1853 504 1943 542
rect 1853 469 1874 504
rect 1906 469 1943 504
rect 1473 155 1561 191
rect 37 129 85 135
rect 65 88 85 129
rect 37 -274 85 88
rect 54 -302 85 -274
rect 37 -310 85 -302
rect 1473 126 1493 155
rect 1522 126 1561 155
rect 1473 -138 1561 126
rect 1473 -167 1492 -138
rect 1521 -167 1561 -138
rect 8 -424 78 -414
rect 1473 -419 1561 -167
rect 1853 -419 1943 469
rect 7 -430 78 -424
rect 6 -459 34 -430
rect 69 -449 78 -430
rect 69 -459 77 -449
rect 6 -816 77 -459
rect 6 -853 18 -816
rect 51 -853 77 -816
rect 6 -860 77 -853
rect 8 -961 82 -948
rect 8 -1010 20 -961
rect 66 -1010 82 -961
rect 8 -1024 82 -1010
rect 9 -1367 82 -1024
rect 9 -1407 18 -1367
rect 53 -1407 82 -1367
rect 9 -1412 82 -1407
<< rmetal3 >>
rect 10 129 37 134
rect 10 88 20 129
rect 10 -274 37 88
rect 10 -302 24 -274
rect 10 -310 37 -302
rect 10 -311 58 -310
use bctr  bctr_0 bitcounter
timestamp 1710559709
transform 1 0 851 0 1 -1106
box -852 -3 1473 541
use bctr  bctr_1
timestamp 1710559709
transform 1 0 856 0 -1 -1129
box -852 -3 1473 541
use bctr  bctr_2
timestamp 1710559709
transform 1 0 847 0 1 6
box -852 -3 1473 541
use bctr  bctr_3
timestamp 1710559709
transform 1 0 854 0 -1 -19
box -852 -3 1473 541
<< end >>
