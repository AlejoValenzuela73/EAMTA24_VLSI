magic
tech sky130A
magscale 1 2
timestamp 1709756558
<< poly >>
rect 72 1026 102 1094
rect 72 408 102 459
<< metal1 >>
rect 28 486 60 1014
rect 114 486 146 1008
use grid  grid_0 grid
timestamp 1678218586
transform 1 0 -9 0 1 266
box -61 -10 259 1053
use sky130_fd_pr__nfet_01v8_NDWVGB  sky130_fd_pr__nfet_01v8_NDWVGB_0
timestamp 1709751578
transform 1 0 87 0 1 435
box -73 -101 73 101
use sky130_fd_pr__pfet_01v8_52N7RA  sky130_fd_pr__pfet_01v8_52N7RA_0
timestamp 1709751578
transform 1 0 87 0 1 1077
box -109 -177 109 177
<< labels >>
rlabel metal1 28 486 60 728 1 in
rlabel metal1 114 486 146 728 1 out
rlabel poly 72 408 102 459 1 clk_2
rlabel poly 72 1026 102 1094 1 clk_1
flabel space -268 1295 -268 1295 0 FreeSans 160 0 0 0 PassGate
<< end >>
