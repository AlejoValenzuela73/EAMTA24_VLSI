magic
tech sky130A
magscale 1 2
timestamp 1710560808
<< nwell >>
rect -1696 1052 -770 1076
rect -78 1074 290 1082
rect -78 1070 306 1074
rect -78 1068 304 1070
rect -1202 1048 -796 1052
rect -1202 1040 -798 1048
rect -662 1040 -282 1042
rect -1202 1008 -282 1040
rect -1202 992 -642 1008
rect -1202 982 -934 992
rect -886 990 -784 992
rect -886 982 -798 990
rect -1202 776 -798 982
rect -1202 652 -958 776
rect -896 732 -798 776
rect -404 732 -54 796
rect -14 732 304 1068
rect -896 728 304 732
rect -896 652 -798 728
rect -1202 560 -798 652
rect -1202 534 -790 560
rect -1202 484 -1120 534
rect -1080 474 -790 534
rect -404 502 -54 728
rect -14 556 304 728
rect -16 520 994 556
rect -16 519 274 520
rect -20 514 274 519
rect -22 508 274 514
rect 420 508 994 520
rect -22 496 218 508
rect -22 490 280 496
rect 512 490 994 508
rect 512 482 698 490
<< poly >>
rect -568 528 -538 538
rect -1052 460 -838 494
rect -916 456 -838 460
<< metal1 >>
rect -662 1040 -282 1042
rect -1100 1008 -282 1040
rect -1100 992 -642 1008
rect -76 998 100 1054
rect -1098 986 -1096 992
rect -1040 896 -866 944
rect -1040 856 -974 896
rect -1072 732 -974 856
rect -1072 672 -1058 732
rect -992 672 -974 732
rect -1072 660 -974 672
rect -1072 440 -1002 660
rect -1064 288 -990 306
rect -1064 222 -1058 288
rect -1006 222 -990 288
rect -1064 164 -990 222
rect -1064 102 -858 164
rect -1014 48 -621 52
rect -1204 10 -621 48
rect -1014 4 -621 10
rect -47 4 135 55
<< via1 >>
rect -1058 672 -992 732
rect -1058 222 -1006 288
<< metal2 >>
rect -1072 732 -848 738
rect -1072 672 -1058 732
rect -992 730 2662 732
rect -992 672 2674 730
rect -1072 668 2674 672
rect -896 666 2674 668
rect -1704 574 -1372 578
rect -1704 504 -1356 574
rect 0 508 70 624
rect -1440 308 -1356 504
rect -104 436 72 508
rect 2610 448 2674 666
rect -1440 306 -1010 308
rect -1440 288 -998 306
rect -1440 236 -1058 288
rect -1436 222 -1058 236
rect -1006 222 -998 288
rect -1436 210 -998 222
use and  and_0 cells
timestamp 1710560808
transform -1 0 -1066 0 1 -6
box -62 0 632 1063
use ffdr3  ffdr3_0 cells
timestamp 1710534732
transform 1 0 322 0 1 2
box -322 -2 2624 1079
use xor  xor_0 cells
timestamp 1710560808
transform 1 0 -662 0 1 0
box -386 -4 652 1074
<< end >>
