magic
tech sky130A
magscale 1 2
timestamp 1710739890
<< nwell >>
rect 16 -848 154 -828
rect 14 -898 156 -848
rect 16 -932 154 -898
rect 4444 -932 4608 -782
rect -10 -1170 4608 -932
rect -10 -1532 4592 -1170
rect 604 -2750 894 -2744
rect 570 -2752 894 -2750
rect 570 -2756 1040 -2752
rect 570 -2760 1674 -2756
rect 2196 -2758 2382 -2752
rect 2070 -2760 2390 -2758
rect 570 -2762 3022 -2760
rect -34 -2764 3022 -2762
rect 3314 -2764 3634 -2762
rect -34 -2766 3634 -2764
rect -34 -2768 3654 -2766
rect -34 -2772 4286 -2768
rect -34 -3349 4590 -2772
rect -34 -3382 4584 -3349
<< nmos >>
rect 812 -2676 842 -2526
rect 908 -2676 938 -2526
rect 1116 -2670 1146 -2370
rect 1212 -2670 1242 -2370
rect 1308 -2670 1338 -2370
rect 1404 -2670 1434 -2370
rect 1870 -2690 1900 -2540
rect 2168 -2636 2198 -2486
rect 2264 -2636 2294 -2486
rect 2694 -2600 2724 -2450
rect 2790 -2600 2820 -2450
rect 3148 -2688 3178 -2538
rect 3432 -2644 3462 -2494
rect 3528 -2644 3558 -2494
rect 3958 -2608 3988 -2458
rect 4054 -2608 4084 -2458
rect 4412 -2696 4442 -2546
<< pmos >>
rect 811 -3128 841 -2828
rect 907 -3128 937 -2828
rect 1116 -3130 1146 -2830
rect 1212 -3130 1242 -2830
rect 1308 -3130 1338 -2830
rect 1404 -3130 1434 -2830
rect 1872 -3156 1902 -2856
rect 2168 -3110 2198 -2810
rect 2264 -3110 2294 -2810
rect 2595 -3138 2625 -2838
rect 2691 -3138 2721 -2838
rect 2787 -3138 2817 -2838
rect 2883 -3138 2913 -2838
rect 3150 -3154 3180 -2854
rect 3432 -3118 3462 -2818
rect 3528 -3118 3558 -2818
rect 3859 -3146 3889 -2846
rect 3955 -3146 3985 -2846
rect 4051 -3146 4081 -2846
rect 4147 -3146 4177 -2846
rect 4414 -3162 4444 -2862
<< ndiff >>
rect 1054 -2382 1116 -2370
rect 750 -2538 812 -2526
rect 750 -2664 762 -2538
rect 796 -2664 812 -2538
rect 750 -2676 812 -2664
rect 842 -2538 908 -2526
rect 842 -2664 858 -2538
rect 892 -2664 908 -2538
rect 842 -2676 908 -2664
rect 938 -2538 1000 -2526
rect 938 -2664 954 -2538
rect 988 -2664 1000 -2538
rect 938 -2676 1000 -2664
rect 1054 -2658 1066 -2382
rect 1100 -2658 1116 -2382
rect 1054 -2670 1116 -2658
rect 1146 -2382 1212 -2370
rect 1146 -2658 1162 -2382
rect 1196 -2658 1212 -2382
rect 1146 -2670 1212 -2658
rect 1242 -2382 1308 -2370
rect 1242 -2658 1258 -2382
rect 1292 -2658 1308 -2382
rect 1242 -2670 1308 -2658
rect 1338 -2382 1404 -2370
rect 1338 -2658 1354 -2382
rect 1388 -2658 1404 -2382
rect 1338 -2670 1404 -2658
rect 1434 -2382 1496 -2370
rect 1434 -2658 1450 -2382
rect 1484 -2658 1496 -2382
rect 2632 -2462 2694 -2450
rect 2106 -2498 2168 -2486
rect 1812 -2552 1870 -2540
rect 1434 -2670 1496 -2658
rect 1812 -2678 1824 -2552
rect 1858 -2678 1870 -2552
rect 1812 -2690 1870 -2678
rect 1900 -2552 1958 -2540
rect 1900 -2678 1912 -2552
rect 1946 -2678 1958 -2552
rect 2106 -2624 2118 -2498
rect 2152 -2624 2168 -2498
rect 2106 -2636 2168 -2624
rect 2198 -2498 2264 -2486
rect 2198 -2624 2214 -2498
rect 2248 -2624 2264 -2498
rect 2198 -2636 2264 -2624
rect 2294 -2498 2356 -2486
rect 2294 -2624 2310 -2498
rect 2344 -2624 2356 -2498
rect 2632 -2588 2644 -2462
rect 2678 -2588 2694 -2462
rect 2632 -2600 2694 -2588
rect 2724 -2462 2790 -2450
rect 2724 -2588 2740 -2462
rect 2774 -2588 2790 -2462
rect 2724 -2600 2790 -2588
rect 2820 -2462 2882 -2450
rect 2820 -2588 2836 -2462
rect 2870 -2588 2882 -2462
rect 3896 -2470 3958 -2458
rect 3370 -2506 3432 -2494
rect 2820 -2600 2882 -2588
rect 3090 -2550 3148 -2538
rect 2294 -2636 2356 -2624
rect 1900 -2690 1958 -2678
rect 3090 -2676 3102 -2550
rect 3136 -2676 3148 -2550
rect 3090 -2688 3148 -2676
rect 3178 -2550 3236 -2538
rect 3178 -2676 3190 -2550
rect 3224 -2676 3236 -2550
rect 3370 -2632 3382 -2506
rect 3416 -2632 3432 -2506
rect 3370 -2644 3432 -2632
rect 3462 -2506 3528 -2494
rect 3462 -2632 3478 -2506
rect 3512 -2632 3528 -2506
rect 3462 -2644 3528 -2632
rect 3558 -2506 3620 -2494
rect 3558 -2632 3574 -2506
rect 3608 -2632 3620 -2506
rect 3896 -2596 3908 -2470
rect 3942 -2596 3958 -2470
rect 3896 -2608 3958 -2596
rect 3988 -2470 4054 -2458
rect 3988 -2596 4004 -2470
rect 4038 -2596 4054 -2470
rect 3988 -2608 4054 -2596
rect 4084 -2470 4146 -2458
rect 4084 -2596 4100 -2470
rect 4134 -2596 4146 -2470
rect 4084 -2608 4146 -2596
rect 4354 -2558 4412 -2546
rect 3558 -2644 3620 -2632
rect 3178 -2688 3236 -2676
rect 4354 -2684 4366 -2558
rect 4400 -2684 4412 -2558
rect 4354 -2696 4412 -2684
rect 4442 -2558 4500 -2546
rect 4442 -2684 4454 -2558
rect 4488 -2684 4500 -2558
rect 4442 -2696 4500 -2684
<< pdiff >>
rect 749 -2840 811 -2828
rect 749 -3116 761 -2840
rect 795 -3116 811 -2840
rect 749 -3128 811 -3116
rect 841 -2840 907 -2828
rect 841 -3116 857 -2840
rect 891 -3116 907 -2840
rect 841 -3128 907 -3116
rect 937 -2840 999 -2828
rect 937 -3116 953 -2840
rect 987 -3116 999 -2840
rect 937 -3128 999 -3116
rect 1054 -2842 1116 -2830
rect 1054 -3118 1066 -2842
rect 1100 -3118 1116 -2842
rect 1054 -3130 1116 -3118
rect 1146 -2842 1212 -2830
rect 1146 -3118 1162 -2842
rect 1196 -3118 1212 -2842
rect 1146 -3130 1212 -3118
rect 1242 -2842 1308 -2830
rect 1242 -3118 1258 -2842
rect 1292 -3118 1308 -2842
rect 1242 -3130 1308 -3118
rect 1338 -2842 1404 -2830
rect 1338 -3118 1354 -2842
rect 1388 -3118 1404 -2842
rect 1338 -3130 1404 -3118
rect 1434 -2842 1496 -2830
rect 1434 -3118 1450 -2842
rect 1484 -3118 1496 -2842
rect 1434 -3130 1496 -3118
rect 2106 -2822 2168 -2810
rect 1814 -2868 1872 -2856
rect 1814 -3144 1826 -2868
rect 1860 -3144 1872 -2868
rect 1814 -3156 1872 -3144
rect 1902 -2868 1960 -2856
rect 1902 -3144 1914 -2868
rect 1948 -3144 1960 -2868
rect 2106 -3098 2118 -2822
rect 2152 -3098 2168 -2822
rect 2106 -3110 2168 -3098
rect 2198 -2822 2264 -2810
rect 2198 -3098 2214 -2822
rect 2248 -3098 2264 -2822
rect 2198 -3110 2264 -3098
rect 2294 -2822 2356 -2810
rect 2294 -3098 2310 -2822
rect 2344 -3098 2356 -2822
rect 2294 -3110 2356 -3098
rect 2533 -2850 2595 -2838
rect 2533 -3126 2545 -2850
rect 2579 -3126 2595 -2850
rect 2533 -3138 2595 -3126
rect 2625 -2850 2691 -2838
rect 2625 -3126 2641 -2850
rect 2675 -3126 2691 -2850
rect 2625 -3138 2691 -3126
rect 2721 -2850 2787 -2838
rect 2721 -3126 2737 -2850
rect 2771 -3126 2787 -2850
rect 2721 -3138 2787 -3126
rect 2817 -2850 2883 -2838
rect 2817 -3126 2833 -2850
rect 2867 -3126 2883 -2850
rect 2817 -3138 2883 -3126
rect 2913 -2850 2975 -2838
rect 2913 -3126 2929 -2850
rect 2963 -3126 2975 -2850
rect 3370 -2830 3432 -2818
rect 2913 -3138 2975 -3126
rect 3092 -2866 3150 -2854
rect 1902 -3156 1960 -3144
rect 3092 -3142 3104 -2866
rect 3138 -3142 3150 -2866
rect 3092 -3154 3150 -3142
rect 3180 -2866 3238 -2854
rect 3180 -3142 3192 -2866
rect 3226 -3142 3238 -2866
rect 3370 -3106 3382 -2830
rect 3416 -3106 3432 -2830
rect 3370 -3118 3432 -3106
rect 3462 -2830 3528 -2818
rect 3462 -3106 3478 -2830
rect 3512 -3106 3528 -2830
rect 3462 -3118 3528 -3106
rect 3558 -2830 3620 -2818
rect 3558 -3106 3574 -2830
rect 3608 -3106 3620 -2830
rect 3558 -3118 3620 -3106
rect 3797 -2858 3859 -2846
rect 3180 -3154 3238 -3142
rect 3797 -3134 3809 -2858
rect 3843 -3134 3859 -2858
rect 3797 -3146 3859 -3134
rect 3889 -2858 3955 -2846
rect 3889 -3134 3905 -2858
rect 3939 -3134 3955 -2858
rect 3889 -3146 3955 -3134
rect 3985 -2858 4051 -2846
rect 3985 -3134 4001 -2858
rect 4035 -3134 4051 -2858
rect 3985 -3146 4051 -3134
rect 4081 -2858 4147 -2846
rect 4081 -3134 4097 -2858
rect 4131 -3134 4147 -2858
rect 4081 -3146 4147 -3134
rect 4177 -2858 4239 -2846
rect 4177 -3134 4193 -2858
rect 4227 -3134 4239 -2858
rect 4177 -3146 4239 -3134
rect 4356 -2874 4414 -2862
rect 4356 -3150 4368 -2874
rect 4402 -3150 4414 -2874
rect 4356 -3162 4414 -3150
rect 4444 -2874 4502 -2862
rect 4444 -3150 4456 -2874
rect 4490 -3150 4502 -2874
rect 4444 -3162 4502 -3150
<< ndiffc >>
rect 762 -2664 796 -2538
rect 858 -2664 892 -2538
rect 954 -2664 988 -2538
rect 1066 -2658 1100 -2382
rect 1162 -2658 1196 -2382
rect 1258 -2658 1292 -2382
rect 1354 -2658 1388 -2382
rect 1450 -2658 1484 -2382
rect 1824 -2678 1858 -2552
rect 1912 -2678 1946 -2552
rect 2118 -2624 2152 -2498
rect 2214 -2624 2248 -2498
rect 2310 -2624 2344 -2498
rect 2644 -2588 2678 -2462
rect 2740 -2588 2774 -2462
rect 2836 -2588 2870 -2462
rect 3102 -2676 3136 -2550
rect 3190 -2676 3224 -2550
rect 3382 -2632 3416 -2506
rect 3478 -2632 3512 -2506
rect 3574 -2632 3608 -2506
rect 3908 -2596 3942 -2470
rect 4004 -2596 4038 -2470
rect 4100 -2596 4134 -2470
rect 4366 -2684 4400 -2558
rect 4454 -2684 4488 -2558
<< pdiffc >>
rect 761 -3116 795 -2840
rect 857 -3116 891 -2840
rect 953 -3116 987 -2840
rect 1066 -3118 1100 -2842
rect 1162 -3118 1196 -2842
rect 1258 -3118 1292 -2842
rect 1354 -3118 1388 -2842
rect 1450 -3118 1484 -2842
rect 1826 -3144 1860 -2868
rect 1914 -3144 1948 -2868
rect 2118 -3098 2152 -2822
rect 2214 -3098 2248 -2822
rect 2310 -3098 2344 -2822
rect 2545 -3126 2579 -2850
rect 2641 -3126 2675 -2850
rect 2737 -3126 2771 -2850
rect 2833 -3126 2867 -2850
rect 2929 -3126 2963 -2850
rect 3104 -3142 3138 -2866
rect 3192 -3142 3226 -2866
rect 3382 -3106 3416 -2830
rect 3478 -3106 3512 -2830
rect 3574 -3106 3608 -2830
rect 3809 -3134 3843 -2858
rect 3905 -3134 3939 -2858
rect 4001 -3134 4035 -2858
rect 4097 -3134 4131 -2858
rect 4193 -3134 4227 -2858
rect 4368 -3150 4402 -2874
rect 4456 -3150 4490 -2874
<< psubdiff >>
rect 21 -2308 45 -2274
rect 245 -2308 269 -2274
rect 333 -2308 357 -2274
rect 557 -2308 581 -2274
rect 737 -2310 761 -2276
rect 961 -2310 985 -2276
rect 1059 -2314 1083 -2280
rect 1283 -2314 1307 -2280
rect 1391 -2316 1415 -2282
rect 1615 -2316 1639 -2282
rect 1765 -2324 1789 -2290
rect 1989 -2324 2013 -2290
rect 2107 -2316 2131 -2282
rect 2331 -2316 2355 -2282
rect 2631 -2324 2655 -2290
rect 2855 -2324 2879 -2290
rect 3043 -2322 3067 -2288
rect 3267 -2322 3291 -2288
rect 3371 -2324 3395 -2290
rect 3595 -2324 3619 -2290
rect 3895 -2332 3919 -2298
rect 4119 -2332 4143 -2298
rect 4307 -2330 4331 -2296
rect 4531 -2330 4555 -2296
<< nsubdiff >>
rect 22 -3256 270 -3255
rect 22 -3290 74 -3256
rect 221 -3290 270 -3256
rect 22 -3291 270 -3290
rect 334 -3256 582 -3255
rect 334 -3290 386 -3256
rect 533 -3290 582 -3256
rect 334 -3291 582 -3290
rect 736 -3258 984 -3257
rect 736 -3292 785 -3258
rect 932 -3292 984 -3258
rect 736 -3293 984 -3292
rect 1058 -3262 1306 -3261
rect 1058 -3296 1107 -3262
rect 1254 -3296 1306 -3262
rect 1058 -3297 1306 -3296
rect 1390 -3264 1638 -3263
rect 1390 -3298 1439 -3264
rect 1586 -3298 1638 -3264
rect 2106 -3264 2354 -3263
rect 1390 -3299 1638 -3298
rect 1764 -3272 2012 -3271
rect 1764 -3306 1813 -3272
rect 1960 -3306 2012 -3272
rect 2106 -3298 2155 -3264
rect 2302 -3298 2354 -3264
rect 3042 -3270 3290 -3269
rect 2106 -3299 2354 -3298
rect 2630 -3272 2878 -3271
rect 1764 -3307 2012 -3306
rect 2630 -3306 2679 -3272
rect 2826 -3306 2878 -3272
rect 3042 -3304 3091 -3270
rect 3238 -3304 3290 -3270
rect 3042 -3305 3290 -3304
rect 3370 -3272 3618 -3271
rect 2630 -3307 2878 -3306
rect 3370 -3306 3419 -3272
rect 3566 -3306 3618 -3272
rect 4306 -3278 4554 -3277
rect 3370 -3307 3618 -3306
rect 3894 -3280 4142 -3279
rect 3894 -3314 3943 -3280
rect 4090 -3314 4142 -3280
rect 4306 -3312 4355 -3278
rect 4502 -3312 4554 -3278
rect 4306 -3313 4554 -3312
rect 3894 -3315 4142 -3314
<< psubdiffcont >>
rect 45 -2308 245 -2274
rect 357 -2308 557 -2274
rect 761 -2310 961 -2276
rect 1083 -2314 1283 -2280
rect 1415 -2316 1615 -2282
rect 1789 -2324 1989 -2290
rect 2131 -2316 2331 -2282
rect 2655 -2324 2855 -2290
rect 3067 -2322 3267 -2288
rect 3395 -2324 3595 -2290
rect 3919 -2332 4119 -2298
rect 4331 -2330 4531 -2296
<< nsubdiffcont >>
rect 74 -3290 221 -3256
rect 386 -3290 533 -3256
rect 785 -3292 932 -3258
rect 1107 -3296 1254 -3262
rect 1439 -3298 1586 -3264
rect 1813 -3306 1960 -3272
rect 2155 -3298 2302 -3264
rect 2679 -3306 2826 -3272
rect 3091 -3304 3238 -3270
rect 3419 -3306 3566 -3272
rect 3943 -3314 4090 -3280
rect 4355 -3312 4502 -3278
<< poly >>
rect 1116 -2370 1146 -2344
rect 1212 -2370 1242 -2344
rect 1308 -2370 1338 -2344
rect 1404 -2370 1434 -2344
rect 756 -2374 824 -2372
rect 900 -2374 940 -2372
rect 734 -2390 940 -2374
rect 734 -2424 774 -2390
rect 808 -2424 940 -2390
rect 734 -2438 940 -2424
rect 756 -2440 824 -2438
rect 900 -2472 940 -2438
rect 906 -2500 940 -2472
rect 812 -2526 842 -2500
rect 908 -2526 938 -2500
rect 2144 -2376 2212 -2358
rect 2144 -2410 2162 -2376
rect 2196 -2410 2212 -2376
rect 2144 -2426 2212 -2410
rect 3506 -2388 3574 -2370
rect 3506 -2422 3524 -2388
rect 3558 -2422 3574 -2388
rect 2168 -2468 2204 -2426
rect 2694 -2450 2724 -2424
rect 2790 -2450 2820 -2424
rect 3506 -2438 3574 -2422
rect 2168 -2486 2198 -2468
rect 2264 -2486 2294 -2460
rect 1870 -2540 1900 -2514
rect 1528 -2612 1596 -2600
rect 1524 -2618 1608 -2612
rect 1524 -2652 1546 -2618
rect 1580 -2652 1608 -2618
rect 812 -2694 842 -2676
rect 908 -2692 938 -2676
rect 1116 -2692 1146 -2670
rect 588 -2718 656 -2710
rect 570 -2728 656 -2718
rect 806 -2726 848 -2694
rect 906 -2710 1146 -2692
rect 570 -2750 604 -2728
rect 588 -2762 604 -2750
rect 638 -2730 656 -2728
rect 768 -2730 848 -2726
rect 638 -2762 848 -2730
rect 588 -2764 848 -2762
rect 588 -2778 656 -2764
rect 718 -2770 848 -2764
rect 806 -2808 848 -2770
rect 902 -2758 1146 -2710
rect 902 -2804 948 -2758
rect 811 -2828 841 -2808
rect 907 -2828 937 -2804
rect 664 -3068 718 -3056
rect 636 -3086 718 -3068
rect 636 -3120 654 -3086
rect 688 -3120 718 -3086
rect 636 -3136 718 -3120
rect 1116 -2830 1146 -2758
rect 1212 -2830 1242 -2670
rect 1308 -2830 1338 -2670
rect 1404 -2688 1434 -2670
rect 1524 -2688 1608 -2652
rect 1402 -2704 1608 -2688
rect 2488 -2518 2604 -2498
rect 2488 -2552 2506 -2518
rect 2540 -2552 2604 -2518
rect 2488 -2612 2604 -2552
rect 3432 -2494 3462 -2468
rect 3528 -2476 3566 -2438
rect 3958 -2458 3988 -2432
rect 4054 -2458 4084 -2432
rect 3528 -2494 3558 -2476
rect 3148 -2538 3178 -2512
rect 2564 -2622 2604 -2612
rect 2694 -2622 2724 -2600
rect 2564 -2624 2724 -2622
rect 1402 -2746 1590 -2704
rect 1870 -2712 1900 -2690
rect 1870 -2732 1902 -2712
rect 1404 -2830 1434 -2746
rect 1716 -2828 1902 -2732
rect 2168 -2810 2198 -2636
rect 2264 -2810 2294 -2636
rect 2564 -2652 2730 -2624
rect 2480 -2722 2630 -2712
rect 2476 -2740 2630 -2722
rect 2476 -2774 2494 -2740
rect 2528 -2770 2630 -2740
rect 2692 -2768 2730 -2652
rect 2790 -2626 2820 -2600
rect 2790 -2656 2920 -2626
rect 2882 -2732 2920 -2656
rect 3752 -2526 3868 -2506
rect 3752 -2560 3770 -2526
rect 3804 -2560 3868 -2526
rect 3752 -2620 3868 -2560
rect 4412 -2546 4442 -2520
rect 3828 -2630 3868 -2620
rect 3958 -2630 3988 -2608
rect 3828 -2632 3988 -2630
rect 3148 -2710 3178 -2688
rect 3148 -2722 3180 -2710
rect 3050 -2726 3180 -2722
rect 2528 -2774 2544 -2770
rect 2476 -2790 2544 -2774
rect 664 -3188 718 -3136
rect 811 -3144 841 -3128
rect 804 -3180 848 -3144
rect 907 -3154 937 -3128
rect 1540 -2850 1608 -2832
rect 1540 -2884 1558 -2850
rect 1592 -2878 1608 -2850
rect 1592 -2884 1616 -2878
rect 1540 -2900 1616 -2884
rect 1116 -3156 1146 -3130
rect 1212 -3158 1242 -3130
rect 1208 -3174 1242 -3158
rect 1308 -3166 1338 -3130
rect 1404 -3160 1434 -3130
rect 1208 -3178 1244 -3174
rect 798 -3188 852 -3180
rect 664 -3204 852 -3188
rect 1202 -3204 1244 -3178
rect 664 -3214 1244 -3204
rect 674 -3228 1244 -3214
rect 798 -3234 1244 -3228
rect 1308 -3214 1346 -3166
rect 1544 -3204 1616 -2900
rect 1718 -3158 1776 -2828
rect 1870 -2838 1902 -2828
rect 1872 -2856 1902 -2838
rect 2588 -2814 2630 -2770
rect 2690 -2812 2818 -2768
rect 2882 -2812 2914 -2732
rect 3048 -2744 3180 -2726
rect 3048 -2778 3066 -2744
rect 3100 -2778 3180 -2744
rect 3048 -2794 3180 -2778
rect 2595 -2838 2625 -2814
rect 2691 -2838 2721 -2812
rect 2786 -2814 2818 -2812
rect 2787 -2838 2817 -2814
rect 2883 -2838 2913 -2812
rect 3148 -2836 3180 -2794
rect 3432 -2818 3462 -2644
rect 3528 -2818 3558 -2644
rect 3828 -2660 3994 -2632
rect 3744 -2730 3894 -2720
rect 3740 -2748 3894 -2730
rect 3740 -2782 3758 -2748
rect 3792 -2778 3894 -2748
rect 3956 -2776 3994 -2660
rect 4054 -2634 4084 -2608
rect 4054 -2664 4184 -2634
rect 4146 -2740 4184 -2664
rect 4412 -2718 4442 -2696
rect 4412 -2730 4444 -2718
rect 4314 -2734 4444 -2730
rect 3792 -2782 3808 -2778
rect 3740 -2798 3808 -2782
rect 2168 -3136 2198 -3110
rect 2264 -3140 2294 -3110
rect 3150 -2854 3180 -2836
rect 1492 -3214 1616 -3204
rect 798 -3236 1240 -3234
rect 1308 -3242 1616 -3214
rect 1702 -3176 1776 -3158
rect 1702 -3210 1720 -3176
rect 1754 -3204 1776 -3176
rect 1872 -3182 1902 -3156
rect 2062 -3172 2130 -3154
rect 1754 -3210 1770 -3204
rect 1702 -3226 1770 -3210
rect 2062 -3206 2080 -3172
rect 2114 -3184 2130 -3172
rect 2262 -3184 2294 -3140
rect 2595 -3164 2625 -3138
rect 2114 -3206 2296 -3184
rect 2062 -3222 2296 -3206
rect 2594 -3210 2626 -3164
rect 2691 -3168 2721 -3138
rect 2787 -3164 2817 -3138
rect 2883 -3156 2913 -3138
rect 3852 -2822 3894 -2778
rect 3954 -2820 4082 -2776
rect 4146 -2820 4178 -2740
rect 4312 -2752 4444 -2734
rect 4312 -2786 4330 -2752
rect 4364 -2786 4444 -2752
rect 4312 -2802 4444 -2786
rect 3859 -2846 3889 -2822
rect 3955 -2846 3985 -2820
rect 4050 -2822 4082 -2820
rect 4051 -2846 4081 -2822
rect 4147 -2846 4177 -2820
rect 4412 -2844 4444 -2802
rect 3432 -3144 3462 -3118
rect 2878 -3210 2914 -3156
rect 3150 -3180 3180 -3154
rect 3422 -3162 3462 -3144
rect 3528 -3148 3558 -3118
rect 4414 -2862 4444 -2844
rect 3326 -3180 3462 -3162
rect 3859 -3172 3889 -3146
rect 2594 -3212 2914 -3210
rect 2594 -3240 2910 -3212
rect 3326 -3214 3344 -3180
rect 3378 -3192 3462 -3180
rect 3378 -3214 3526 -3192
rect 3326 -3230 3526 -3214
rect 3858 -3218 3890 -3172
rect 3955 -3176 3985 -3146
rect 4051 -3172 4081 -3146
rect 4147 -3164 4177 -3146
rect 4142 -3218 4178 -3164
rect 4414 -3188 4444 -3162
rect 3858 -3220 4178 -3218
rect 1308 -3244 1578 -3242
rect 3858 -3248 4174 -3220
<< polycont >>
rect 774 -2424 808 -2390
rect 2162 -2410 2196 -2376
rect 3524 -2422 3558 -2388
rect 1546 -2652 1580 -2618
rect 604 -2762 638 -2728
rect 654 -3120 688 -3086
rect 2506 -2552 2540 -2518
rect 2494 -2774 2528 -2740
rect 3770 -2560 3804 -2526
rect 1558 -2884 1592 -2850
rect 3066 -2778 3100 -2744
rect 3758 -2782 3792 -2748
rect 1720 -3210 1754 -3176
rect 2080 -3206 2114 -3172
rect 4330 -2786 4364 -2752
rect 3344 -3214 3378 -3180
<< locali >>
rect 762 -2390 820 -2372
rect 762 -2424 774 -2390
rect 808 -2424 820 -2390
rect 762 -2440 820 -2424
rect 1066 -2382 1100 -2366
rect 762 -2538 796 -2522
rect 762 -2680 796 -2664
rect 858 -2538 892 -2522
rect 858 -2680 892 -2664
rect 954 -2538 988 -2522
rect 954 -2680 988 -2664
rect 1066 -2674 1100 -2658
rect 1162 -2382 1196 -2366
rect 1162 -2674 1196 -2658
rect 1258 -2382 1292 -2366
rect 1258 -2674 1292 -2658
rect 1354 -2382 1388 -2366
rect 1354 -2674 1388 -2658
rect 1450 -2382 1484 -2366
rect 2150 -2376 2208 -2358
rect 2150 -2410 2162 -2376
rect 2196 -2410 2208 -2376
rect 2150 -2426 2208 -2410
rect 3512 -2388 3570 -2370
rect 3512 -2422 3524 -2388
rect 3558 -2422 3570 -2388
rect 3512 -2438 3570 -2422
rect 2644 -2462 2678 -2446
rect 2118 -2498 2152 -2482
rect 1824 -2552 1858 -2536
rect 1450 -2674 1484 -2658
rect 1534 -2618 1592 -2600
rect 1534 -2652 1546 -2618
rect 1580 -2652 1592 -2618
rect 1534 -2668 1592 -2652
rect 1824 -2694 1858 -2678
rect 1912 -2552 1946 -2536
rect 2118 -2640 2152 -2624
rect 2214 -2498 2248 -2482
rect 2214 -2640 2248 -2624
rect 2310 -2498 2344 -2482
rect 2494 -2518 2552 -2500
rect 2494 -2552 2506 -2518
rect 2540 -2552 2552 -2518
rect 2494 -2568 2552 -2552
rect 2644 -2604 2678 -2588
rect 2740 -2462 2774 -2446
rect 2740 -2604 2774 -2588
rect 2836 -2462 2870 -2446
rect 3908 -2470 3942 -2454
rect 3382 -2506 3416 -2490
rect 2836 -2604 2870 -2588
rect 3102 -2550 3136 -2534
rect 2310 -2640 2344 -2624
rect 1912 -2694 1946 -2678
rect 3102 -2692 3136 -2676
rect 3190 -2550 3224 -2534
rect 3382 -2648 3416 -2632
rect 3478 -2506 3512 -2490
rect 3478 -2648 3512 -2632
rect 3574 -2506 3608 -2490
rect 3758 -2526 3816 -2508
rect 3758 -2560 3770 -2526
rect 3804 -2560 3816 -2526
rect 3758 -2576 3816 -2560
rect 3908 -2612 3942 -2596
rect 4004 -2470 4038 -2454
rect 4004 -2612 4038 -2596
rect 4100 -2470 4134 -2454
rect 4100 -2612 4134 -2596
rect 4366 -2558 4400 -2542
rect 3574 -2648 3608 -2632
rect 3190 -2692 3224 -2676
rect 4366 -2700 4400 -2684
rect 4454 -2558 4488 -2542
rect 4454 -2700 4488 -2684
rect 592 -2728 650 -2710
rect 592 -2762 604 -2728
rect 638 -2762 650 -2728
rect 592 -2778 650 -2762
rect 2482 -2740 2540 -2722
rect 2482 -2774 2494 -2740
rect 2528 -2774 2540 -2740
rect 2482 -2790 2540 -2774
rect 3054 -2744 3112 -2726
rect 3054 -2778 3066 -2744
rect 3100 -2778 3112 -2744
rect 3054 -2794 3112 -2778
rect 3746 -2748 3804 -2730
rect 3746 -2782 3758 -2748
rect 3792 -2782 3804 -2748
rect 3746 -2798 3804 -2782
rect 4318 -2752 4376 -2734
rect 4318 -2786 4330 -2752
rect 4364 -2786 4376 -2752
rect 4318 -2802 4376 -2786
rect 2118 -2822 2152 -2806
rect 761 -2840 795 -2824
rect 642 -3086 700 -3068
rect 642 -3120 654 -3086
rect 688 -3120 700 -3086
rect 642 -3136 700 -3120
rect 761 -3132 795 -3116
rect 857 -2840 891 -2824
rect 857 -3132 891 -3116
rect 953 -2840 987 -2824
rect 953 -3132 987 -3116
rect 1066 -2842 1100 -2826
rect 1066 -3134 1100 -3118
rect 1162 -2842 1196 -2826
rect 1162 -3134 1196 -3118
rect 1258 -2842 1292 -2826
rect 1258 -3134 1292 -3118
rect 1354 -2842 1388 -2826
rect 1354 -3134 1388 -3118
rect 1450 -2842 1484 -2826
rect 1546 -2850 1604 -2832
rect 1546 -2884 1558 -2850
rect 1592 -2884 1604 -2850
rect 1546 -2900 1604 -2884
rect 1826 -2868 1860 -2852
rect 1450 -3134 1484 -3118
rect 1708 -3176 1766 -3158
rect 1826 -3160 1860 -3144
rect 1914 -2868 1948 -2852
rect 2118 -3114 2152 -3098
rect 2214 -2822 2248 -2806
rect 2214 -3114 2248 -3098
rect 2310 -2822 2344 -2806
rect 3382 -2830 3416 -2814
rect 2310 -3114 2344 -3098
rect 2545 -2850 2579 -2834
rect 2545 -3142 2579 -3126
rect 2641 -2850 2675 -2834
rect 2641 -3142 2675 -3126
rect 2737 -2850 2771 -2834
rect 2737 -3142 2771 -3126
rect 2833 -2850 2867 -2834
rect 2833 -3142 2867 -3126
rect 2929 -2850 2963 -2834
rect 2929 -3142 2963 -3126
rect 3104 -2866 3138 -2850
rect 1914 -3160 1948 -3144
rect 1708 -3210 1720 -3176
rect 1754 -3210 1766 -3176
rect 1708 -3226 1766 -3210
rect 2068 -3172 2126 -3154
rect 3104 -3158 3138 -3142
rect 3192 -2866 3226 -2850
rect 3382 -3122 3416 -3106
rect 3478 -2830 3512 -2814
rect 3478 -3122 3512 -3106
rect 3574 -2830 3608 -2814
rect 3574 -3122 3608 -3106
rect 3809 -2858 3843 -2842
rect 3192 -3158 3226 -3142
rect 3809 -3150 3843 -3134
rect 3905 -2858 3939 -2842
rect 3905 -3150 3939 -3134
rect 4001 -2858 4035 -2842
rect 4001 -3150 4035 -3134
rect 4097 -2858 4131 -2842
rect 4097 -3150 4131 -3134
rect 4193 -2858 4227 -2842
rect 4193 -3150 4227 -3134
rect 4368 -2874 4402 -2858
rect 2068 -3206 2080 -3172
rect 2114 -3206 2126 -3172
rect 2068 -3222 2126 -3206
rect 3332 -3180 3390 -3162
rect 4368 -3166 4402 -3150
rect 4456 -2874 4490 -2858
rect 4456 -3166 4490 -3150
rect 3332 -3214 3344 -3180
rect 3378 -3214 3390 -3180
rect 3332 -3230 3390 -3214
rect 13 -3252 279 -3248
rect 13 -3295 18 -3252
rect 273 -3295 279 -3252
rect 13 -3298 279 -3295
rect 325 -3252 591 -3248
rect 325 -3295 330 -3252
rect 585 -3295 591 -3252
rect 325 -3298 591 -3295
rect 727 -3254 993 -3250
rect 727 -3297 733 -3254
rect 988 -3297 993 -3254
rect 727 -3300 993 -3297
rect 1049 -3258 1315 -3254
rect 1049 -3301 1055 -3258
rect 1310 -3301 1315 -3258
rect 1049 -3304 1315 -3301
rect 1381 -3260 1647 -3256
rect 1381 -3303 1387 -3260
rect 1642 -3303 1647 -3260
rect 2097 -3260 2363 -3256
rect 1381 -3306 1647 -3303
rect 1755 -3268 2021 -3264
rect 1755 -3311 1761 -3268
rect 2016 -3311 2021 -3268
rect 2097 -3303 2103 -3260
rect 2358 -3303 2363 -3260
rect 2097 -3306 2363 -3303
rect 2621 -3268 2887 -3264
rect 1755 -3314 2021 -3311
rect 2621 -3311 2627 -3268
rect 2882 -3311 2887 -3268
rect 2621 -3314 2887 -3311
rect 3033 -3266 3299 -3262
rect 3033 -3309 3039 -3266
rect 3294 -3309 3299 -3266
rect 3033 -3312 3299 -3309
rect 3361 -3268 3627 -3264
rect 3361 -3311 3367 -3268
rect 3622 -3311 3627 -3268
rect 3361 -3314 3627 -3311
rect 3885 -3276 4151 -3272
rect 3885 -3319 3891 -3276
rect 4146 -3319 4151 -3276
rect 3885 -3322 4151 -3319
rect 4297 -3274 4563 -3270
rect 4297 -3317 4303 -3274
rect 4558 -3317 4563 -3274
rect 4297 -3320 4563 -3317
<< viali >>
rect 17 -2274 272 -2270
rect 17 -2308 45 -2274
rect 45 -2308 245 -2274
rect 245 -2308 272 -2274
rect 17 -2313 272 -2308
rect 329 -2274 584 -2270
rect 329 -2308 357 -2274
rect 357 -2308 557 -2274
rect 557 -2308 584 -2274
rect 329 -2313 584 -2308
rect 734 -2276 989 -2272
rect 734 -2310 761 -2276
rect 761 -2310 961 -2276
rect 961 -2310 989 -2276
rect 734 -2315 989 -2310
rect 1056 -2280 1311 -2276
rect 1056 -2314 1083 -2280
rect 1083 -2314 1283 -2280
rect 1283 -2314 1311 -2280
rect 1056 -2319 1311 -2314
rect 1388 -2282 1643 -2278
rect 1388 -2316 1415 -2282
rect 1415 -2316 1615 -2282
rect 1615 -2316 1643 -2282
rect 2104 -2282 2359 -2278
rect 1388 -2321 1643 -2316
rect 1762 -2290 2017 -2286
rect 1762 -2324 1789 -2290
rect 1789 -2324 1989 -2290
rect 1989 -2324 2017 -2290
rect 2104 -2316 2131 -2282
rect 2131 -2316 2331 -2282
rect 2331 -2316 2359 -2282
rect 2104 -2321 2359 -2316
rect 2628 -2290 2883 -2286
rect 1762 -2329 2017 -2324
rect 2628 -2324 2655 -2290
rect 2655 -2324 2855 -2290
rect 2855 -2324 2883 -2290
rect 2628 -2329 2883 -2324
rect 3040 -2288 3295 -2284
rect 3040 -2322 3067 -2288
rect 3067 -2322 3267 -2288
rect 3267 -2322 3295 -2288
rect 3040 -2327 3295 -2322
rect 3368 -2290 3623 -2286
rect 3368 -2324 3395 -2290
rect 3395 -2324 3595 -2290
rect 3595 -2324 3623 -2290
rect 3368 -2329 3623 -2324
rect 3892 -2298 4147 -2294
rect 3892 -2332 3919 -2298
rect 3919 -2332 4119 -2298
rect 4119 -2332 4147 -2298
rect 3892 -2337 4147 -2332
rect 4304 -2296 4559 -2292
rect 4304 -2330 4331 -2296
rect 4331 -2330 4531 -2296
rect 4531 -2330 4559 -2296
rect 4304 -2335 4559 -2330
rect 774 -2424 808 -2390
rect 762 -2664 796 -2538
rect 858 -2664 892 -2538
rect 954 -2664 988 -2538
rect 1066 -2658 1100 -2382
rect 1162 -2658 1196 -2382
rect 1258 -2658 1292 -2382
rect 1354 -2658 1388 -2382
rect 1450 -2658 1484 -2382
rect 2162 -2410 2196 -2376
rect 3524 -2422 3558 -2388
rect 1546 -2652 1580 -2618
rect 1824 -2678 1858 -2552
rect 1912 -2678 1946 -2552
rect 2118 -2624 2152 -2498
rect 2214 -2624 2248 -2498
rect 2310 -2624 2344 -2498
rect 2506 -2552 2540 -2518
rect 2644 -2588 2678 -2462
rect 2740 -2588 2774 -2462
rect 2836 -2588 2870 -2462
rect 3102 -2676 3136 -2550
rect 3190 -2676 3224 -2550
rect 3382 -2632 3416 -2506
rect 3478 -2632 3512 -2506
rect 3574 -2632 3608 -2506
rect 3770 -2560 3804 -2526
rect 3908 -2596 3942 -2470
rect 4004 -2596 4038 -2470
rect 4100 -2596 4134 -2470
rect 4366 -2684 4400 -2558
rect 4454 -2684 4488 -2558
rect 604 -2762 638 -2728
rect 2494 -2774 2528 -2740
rect 3066 -2778 3100 -2744
rect 3758 -2782 3792 -2748
rect 4330 -2786 4364 -2752
rect 654 -3120 688 -3086
rect 761 -3116 795 -2840
rect 857 -3116 891 -2840
rect 953 -3116 987 -2840
rect 1066 -3118 1100 -2842
rect 1162 -3118 1196 -2842
rect 1258 -3118 1292 -2842
rect 1354 -3118 1388 -2842
rect 1450 -3118 1484 -2842
rect 1558 -2884 1592 -2850
rect 1826 -3144 1860 -2868
rect 1914 -3144 1948 -2868
rect 2118 -3098 2152 -2822
rect 2214 -3098 2248 -2822
rect 2310 -3098 2344 -2822
rect 2545 -3126 2579 -2850
rect 2641 -3126 2675 -2850
rect 2737 -3126 2771 -2850
rect 2833 -3126 2867 -2850
rect 2929 -3126 2963 -2850
rect 3104 -3142 3138 -2866
rect 1720 -3210 1754 -3176
rect 3192 -3142 3226 -2866
rect 3382 -3106 3416 -2830
rect 3478 -3106 3512 -2830
rect 3574 -3106 3608 -2830
rect 3809 -3134 3843 -2858
rect 3905 -3134 3939 -2858
rect 4001 -3134 4035 -2858
rect 4097 -3134 4131 -2858
rect 4193 -3134 4227 -2858
rect 4368 -3150 4402 -2874
rect 2080 -3206 2114 -3172
rect 4456 -3150 4490 -2874
rect 3344 -3214 3378 -3180
rect 18 -3256 273 -3252
rect 18 -3290 74 -3256
rect 74 -3290 221 -3256
rect 221 -3290 273 -3256
rect 18 -3295 273 -3290
rect 330 -3256 585 -3252
rect 330 -3290 386 -3256
rect 386 -3290 533 -3256
rect 533 -3290 585 -3256
rect 330 -3295 585 -3290
rect 733 -3258 988 -3254
rect 733 -3292 785 -3258
rect 785 -3292 932 -3258
rect 932 -3292 988 -3258
rect 733 -3297 988 -3292
rect 1055 -3262 1310 -3258
rect 1055 -3296 1107 -3262
rect 1107 -3296 1254 -3262
rect 1254 -3296 1310 -3262
rect 1055 -3301 1310 -3296
rect 1387 -3264 1642 -3260
rect 1387 -3298 1439 -3264
rect 1439 -3298 1586 -3264
rect 1586 -3298 1642 -3264
rect 1387 -3303 1642 -3298
rect 1761 -3272 2016 -3268
rect 1761 -3306 1813 -3272
rect 1813 -3306 1960 -3272
rect 1960 -3306 2016 -3272
rect 1761 -3311 2016 -3306
rect 2103 -3264 2358 -3260
rect 2103 -3298 2155 -3264
rect 2155 -3298 2302 -3264
rect 2302 -3298 2358 -3264
rect 2103 -3303 2358 -3298
rect 2627 -3272 2882 -3268
rect 2627 -3306 2679 -3272
rect 2679 -3306 2826 -3272
rect 2826 -3306 2882 -3272
rect 2627 -3311 2882 -3306
rect 3039 -3270 3294 -3266
rect 3039 -3304 3091 -3270
rect 3091 -3304 3238 -3270
rect 3238 -3304 3294 -3270
rect 3039 -3309 3294 -3304
rect 3367 -3272 3622 -3268
rect 3367 -3306 3419 -3272
rect 3419 -3306 3566 -3272
rect 3566 -3306 3622 -3272
rect 3367 -3311 3622 -3306
rect 3891 -3280 4146 -3276
rect 3891 -3314 3943 -3280
rect 3943 -3314 4090 -3280
rect 4090 -3314 4146 -3280
rect 3891 -3319 4146 -3314
rect 4303 -3278 4558 -3274
rect 4303 -3312 4355 -3278
rect 4355 -3312 4502 -3278
rect 4502 -3312 4558 -3278
rect 4303 -3317 4558 -3312
<< metal1 >>
rect -28 1110 4622 1120
rect -28 1088 4652 1110
rect -28 1032 1512 1088
rect 1580 1032 4652 1088
rect -28 1020 4652 1032
rect 4 258 170 288
rect 4 176 40 258
rect 130 176 170 258
rect 4 128 170 176
rect 40 52 382 58
rect 2 48 4644 52
rect -62 42 4644 48
rect -62 -62 2100 42
rect 2184 -62 4644 42
rect -62 -84 4644 -62
rect -62 -102 138 -84
rect 42 -856 184 -812
rect 42 -922 66 -856
rect 142 -922 184 -856
rect 42 -974 184 -922
rect 38 -1038 4598 -1036
rect 38 -1090 4652 -1038
rect 38 -1146 1510 -1090
rect 1586 -1146 4652 -1090
rect 38 -1214 4652 -1146
rect 38 -1218 3886 -1214
rect 4196 -1218 4652 -1214
rect 4556 -1240 4652 -1218
rect 16 -1922 164 -1868
rect 16 -2020 40 -1922
rect 132 -2020 164 -1922
rect 16 -2058 164 -2020
rect -62 -2144 24 -2142
rect -62 -2166 598 -2144
rect 744 -2166 1018 -2146
rect 1026 -2166 4622 -2164
rect -62 -2206 4632 -2166
rect -62 -2270 2094 -2206
rect -62 -2292 17 -2270
rect -22 -2313 17 -2292
rect 272 -2313 329 -2270
rect 584 -2272 2094 -2270
rect 584 -2313 734 -2272
rect -22 -2314 734 -2313
rect -20 -2315 734 -2314
rect 989 -2276 2094 -2272
rect 989 -2315 1056 -2276
rect -20 -2319 1056 -2315
rect 1311 -2278 2094 -2276
rect 2184 -2278 4632 -2206
rect 1311 -2319 1388 -2278
rect -20 -2321 1388 -2319
rect 1643 -2282 2094 -2278
rect 1643 -2286 2104 -2282
rect 1643 -2321 1762 -2286
rect -20 -2322 1762 -2321
rect -20 -2324 696 -2322
rect 620 -2390 826 -2372
rect 620 -2424 774 -2390
rect 808 -2424 826 -2390
rect 620 -2434 826 -2424
rect 620 -2492 694 -2434
rect 762 -2440 820 -2434
rect 620 -2558 626 -2492
rect 678 -2558 694 -2492
rect 620 -2576 694 -2558
rect 740 -2538 806 -2490
rect 856 -2526 908 -2322
rect 1044 -2324 1762 -2322
rect 1044 -2325 1323 -2324
rect 1376 -2325 1762 -2324
rect 1060 -2370 1102 -2325
rect 1376 -2327 1655 -2325
rect 1446 -2370 1486 -2327
rect 1742 -2329 1762 -2325
rect 2017 -2321 2104 -2286
rect 2359 -2284 4632 -2278
rect 2359 -2286 3040 -2284
rect 2359 -2321 2628 -2286
rect 2017 -2329 2628 -2321
rect 2883 -2327 3040 -2286
rect 3295 -2286 4632 -2284
rect 3295 -2327 3368 -2286
rect 2883 -2329 3368 -2327
rect 3623 -2292 4632 -2286
rect 3623 -2294 4304 -2292
rect 3623 -2329 3892 -2294
rect 1742 -2330 3892 -2329
rect 1750 -2335 2029 -2330
rect 2616 -2335 2895 -2330
rect 3028 -2333 3307 -2330
rect 1060 -2382 1106 -2370
rect 740 -2616 762 -2538
rect 796 -2616 806 -2538
rect 740 -2668 744 -2616
rect 802 -2668 806 -2616
rect 582 -2710 670 -2706
rect 582 -2712 682 -2710
rect 582 -2782 588 -2712
rect 664 -2782 682 -2712
rect 582 -2788 682 -2782
rect 612 -2930 682 -2788
rect 740 -2840 806 -2668
rect 852 -2528 908 -2526
rect 852 -2538 898 -2528
rect 852 -2664 858 -2538
rect 892 -2664 898 -2538
rect 852 -2676 898 -2664
rect 944 -2538 1002 -2498
rect 944 -2664 954 -2538
rect 988 -2664 1002 -2538
rect 944 -2722 1002 -2664
rect 1060 -2658 1066 -2382
rect 1100 -2658 1106 -2382
rect 1060 -2670 1106 -2658
rect 1156 -2382 1202 -2370
rect 1156 -2658 1162 -2382
rect 1196 -2658 1202 -2382
rect 1156 -2670 1202 -2658
rect 1252 -2382 1298 -2370
rect 1252 -2658 1258 -2382
rect 1292 -2658 1298 -2382
rect 1252 -2670 1298 -2658
rect 1348 -2382 1394 -2370
rect 1348 -2658 1354 -2382
rect 1388 -2658 1394 -2382
rect 1348 -2670 1394 -2658
rect 1444 -2382 1490 -2370
rect 1444 -2658 1450 -2382
rect 1484 -2658 1490 -2382
rect 1814 -2552 1866 -2335
rect 2150 -2360 2208 -2358
rect 2144 -2364 2214 -2360
rect 1910 -2368 2214 -2364
rect 1910 -2392 2154 -2368
rect 1444 -2670 1490 -2658
rect 1534 -2610 1592 -2600
rect 1534 -2662 1536 -2610
rect 1588 -2662 1592 -2610
rect 1534 -2668 1592 -2662
rect 1254 -2674 1298 -2670
rect 1254 -2704 1296 -2674
rect 1814 -2678 1824 -2552
rect 1858 -2678 1866 -2552
rect 1814 -2690 1866 -2678
rect 1906 -2420 2154 -2392
rect 2206 -2420 2214 -2368
rect 1906 -2426 2214 -2420
rect 1906 -2440 2208 -2426
rect 1906 -2548 1958 -2440
rect 2620 -2450 2678 -2335
rect 2620 -2462 2684 -2450
rect 2620 -2466 2644 -2462
rect 2406 -2486 2446 -2480
rect 2014 -2498 2158 -2486
rect 1906 -2552 1952 -2548
rect 1906 -2678 1912 -2552
rect 1946 -2622 1952 -2552
rect 1946 -2678 1966 -2622
rect 1906 -2690 1966 -2678
rect 1254 -2714 1674 -2704
rect 926 -2746 1024 -2722
rect 1254 -2742 1586 -2714
rect 926 -2798 948 -2746
rect 1000 -2798 1024 -2746
rect 1348 -2766 1586 -2742
rect 1638 -2766 1674 -2714
rect 926 -2808 1024 -2798
rect 1060 -2802 1298 -2774
rect 740 -2860 761 -2840
rect 612 -2942 710 -2930
rect 612 -3002 626 -2942
rect 692 -3002 710 -2942
rect 612 -3086 710 -3002
rect 612 -3120 654 -3086
rect 688 -3120 710 -3086
rect 612 -3126 710 -3120
rect 642 -3136 710 -3126
rect 755 -3116 761 -2860
rect 795 -2860 806 -2840
rect 851 -2840 897 -2828
rect 795 -3116 801 -2860
rect 755 -3128 801 -3116
rect 851 -3116 857 -2840
rect 891 -3116 897 -2840
rect 944 -2840 1002 -2808
rect 944 -2866 953 -2840
rect 851 -3122 897 -3116
rect 947 -3116 953 -2866
rect 987 -2866 1002 -2840
rect 1060 -2842 1106 -2802
rect 987 -3116 993 -2866
rect 947 -3118 993 -3116
rect 1060 -3118 1066 -2842
rect 1100 -3118 1106 -2842
rect 851 -3128 898 -3122
rect 947 -3128 994 -3118
rect 644 -3166 710 -3136
rect 644 -3214 818 -3166
rect 214 -3246 264 -3222
rect 340 -3246 392 -3222
rect 6 -3248 285 -3246
rect 318 -3248 597 -3246
rect 858 -3248 898 -3128
rect 950 -3156 994 -3128
rect 1060 -3130 1106 -3118
rect 1156 -2842 1202 -2830
rect 1156 -3118 1162 -2842
rect 1196 -3118 1202 -2842
rect 950 -3214 992 -3156
rect 6 -3252 597 -3248
rect 6 -3295 18 -3252
rect 273 -3295 330 -3252
rect 585 -3262 597 -3252
rect 721 -3254 1000 -3248
rect 1156 -3252 1202 -3118
rect 1252 -2842 1298 -2802
rect 1252 -3118 1258 -2842
rect 1292 -3118 1298 -2842
rect 1252 -3192 1298 -3118
rect 1348 -2776 1674 -2766
rect 1348 -2842 1394 -2776
rect 1348 -3118 1354 -2842
rect 1388 -3118 1394 -2842
rect 1348 -3130 1394 -3118
rect 1444 -2842 1490 -2830
rect 1444 -3118 1450 -2842
rect 1484 -3118 1490 -2842
rect 1546 -2838 1604 -2832
rect 1546 -2890 1550 -2838
rect 1602 -2890 1604 -2838
rect 1914 -2856 1966 -2690
rect 2014 -2624 2118 -2498
rect 2152 -2624 2158 -2498
rect 2014 -2636 2158 -2624
rect 2208 -2498 2254 -2486
rect 2208 -2624 2214 -2498
rect 2248 -2624 2254 -2498
rect 2014 -2642 2156 -2636
rect 2014 -2776 2086 -2642
rect 2208 -2678 2254 -2624
rect 2302 -2498 2446 -2486
rect 2302 -2624 2310 -2498
rect 2344 -2624 2446 -2498
rect 2494 -2502 2552 -2500
rect 2490 -2510 2556 -2502
rect 2490 -2562 2496 -2510
rect 2548 -2562 2556 -2510
rect 2490 -2568 2556 -2562
rect 2638 -2588 2644 -2466
rect 2678 -2588 2684 -2462
rect 2734 -2462 2780 -2450
rect 2828 -2458 2894 -2335
rect 2734 -2580 2740 -2462
rect 2638 -2600 2684 -2588
rect 2730 -2588 2740 -2580
rect 2774 -2588 2780 -2462
rect 2302 -2634 2446 -2624
rect 2304 -2636 2350 -2634
rect 2208 -2692 2316 -2678
rect 2208 -2748 2228 -2692
rect 2290 -2748 2316 -2692
rect 2208 -2768 2316 -2748
rect 2014 -2822 2078 -2776
rect 1546 -2900 1604 -2890
rect 1820 -2868 1866 -2856
rect 1820 -2942 1826 -2868
rect 1444 -3164 1490 -3118
rect 1814 -3144 1826 -2942
rect 1860 -3144 1866 -2868
rect 1708 -3164 1766 -3158
rect 1436 -3166 1490 -3164
rect 1436 -3192 1488 -3166
rect 1252 -3220 1488 -3192
rect 1706 -3172 1772 -3164
rect 1706 -3224 1712 -3172
rect 1764 -3224 1772 -3172
rect 1706 -3230 1772 -3224
rect 721 -3262 733 -3254
rect 585 -3295 733 -3262
rect 6 -3297 733 -3295
rect 988 -3262 1000 -3254
rect 1036 -3254 1492 -3252
rect 1036 -3258 1654 -3254
rect 1036 -3262 1055 -3258
rect 988 -3297 1055 -3262
rect 6 -3301 1055 -3297
rect 1310 -3260 1654 -3258
rect 1310 -3301 1387 -3260
rect 1642 -3268 1654 -3260
rect 1814 -3262 1866 -3144
rect 1908 -2868 1966 -2856
rect 1908 -3144 1914 -2868
rect 1948 -3002 1966 -2868
rect 2010 -2830 2078 -2822
rect 2010 -2882 2020 -2830
rect 2072 -2882 2078 -2830
rect 2010 -2888 2078 -2882
rect 2106 -2810 2156 -2804
rect 2106 -2822 2158 -2810
rect 2106 -2892 2118 -2822
rect 1948 -3144 1954 -3002
rect 2112 -3040 2118 -2892
rect 2088 -3048 2118 -3040
rect 2088 -3100 2098 -3048
rect 2152 -3098 2158 -2822
rect 2150 -3100 2158 -3098
rect 2088 -3106 2158 -3100
rect 2112 -3110 2158 -3106
rect 2208 -2822 2254 -2768
rect 2208 -3098 2214 -2822
rect 2248 -3098 2254 -2822
rect 2208 -3110 2254 -3098
rect 2304 -2820 2350 -2810
rect 2304 -2822 2378 -2820
rect 2304 -3098 2310 -2822
rect 2344 -2828 2378 -2822
rect 2370 -2880 2378 -2828
rect 2344 -2886 2378 -2880
rect 2406 -2884 2446 -2634
rect 2730 -2690 2780 -2588
rect 2830 -2462 2876 -2458
rect 2830 -2588 2836 -2462
rect 2870 -2588 2876 -2462
rect 2830 -2600 2876 -2588
rect 3092 -2550 3144 -2333
rect 3354 -2340 3646 -2330
rect 3818 -2337 3892 -2330
rect 4147 -2330 4304 -2294
rect 4147 -2337 4201 -2330
rect 4292 -2335 4304 -2330
rect 4559 -2310 4632 -2292
rect 4559 -2316 4620 -2310
rect 4559 -2335 4571 -2316
rect 3880 -2343 4159 -2337
rect 4292 -2341 4571 -2335
rect 3512 -2372 3570 -2370
rect 3506 -2380 3576 -2372
rect 3506 -2432 3516 -2380
rect 3568 -2432 3576 -2380
rect 3506 -2438 3576 -2432
rect 3884 -2458 3942 -2343
rect 3884 -2470 3948 -2458
rect 3884 -2474 3908 -2470
rect 3670 -2494 3710 -2488
rect 3278 -2506 3422 -2494
rect 3092 -2676 3102 -2550
rect 3136 -2676 3144 -2550
rect 3092 -2688 3144 -2676
rect 3184 -2550 3230 -2538
rect 3184 -2676 3190 -2550
rect 3224 -2620 3230 -2550
rect 3224 -2676 3244 -2620
rect 3184 -2688 3244 -2676
rect 2730 -2710 2784 -2690
rect 2728 -2714 3016 -2710
rect 2728 -2716 3018 -2714
rect 2474 -2730 2548 -2718
rect 2474 -2782 2480 -2730
rect 2532 -2782 2548 -2730
rect 2728 -2722 3106 -2716
rect 2728 -2728 3112 -2722
rect 2728 -2764 2982 -2728
rect 2474 -2790 2548 -2782
rect 2730 -2796 2784 -2764
rect 2930 -2780 2982 -2764
rect 3034 -2744 3112 -2728
rect 3034 -2778 3066 -2744
rect 3100 -2778 3112 -2744
rect 3034 -2780 3112 -2778
rect 2930 -2796 3112 -2780
rect 2539 -2850 2585 -2838
rect 2344 -3098 2350 -2886
rect 2406 -3038 2454 -2884
rect 2304 -3110 2350 -3098
rect 2382 -3046 2454 -3038
rect 2382 -3098 2392 -3046
rect 2444 -3098 2454 -3046
rect 2382 -3104 2454 -3098
rect 2539 -3102 2545 -2850
rect 1908 -3156 1954 -3144
rect 2528 -3126 2545 -3102
rect 2579 -3102 2585 -2850
rect 2635 -2850 2681 -2838
rect 2730 -2848 2780 -2796
rect 2579 -3126 2586 -3102
rect 2068 -3156 2126 -3154
rect 2060 -3164 2130 -3156
rect 2060 -3216 2070 -3164
rect 2122 -3216 2130 -3164
rect 2528 -3172 2586 -3126
rect 2635 -3126 2641 -2850
rect 2675 -3126 2681 -2850
rect 2635 -3136 2681 -3126
rect 2731 -2850 2777 -2848
rect 2731 -3126 2737 -2850
rect 2771 -3126 2777 -2850
rect 2060 -3222 2130 -3216
rect 2091 -3260 2370 -3254
rect 2530 -3260 2582 -3172
rect 2634 -3190 2682 -3136
rect 2731 -3138 2777 -3126
rect 2827 -2850 2873 -2838
rect 2827 -3126 2833 -2850
rect 2867 -3126 2873 -2850
rect 2827 -3138 2873 -3126
rect 2923 -2850 2969 -2838
rect 2923 -3126 2929 -2850
rect 2963 -3126 2969 -2850
rect 3192 -2854 3244 -2688
rect 3278 -2632 3382 -2506
rect 3416 -2632 3422 -2506
rect 3278 -2644 3422 -2632
rect 3472 -2506 3518 -2494
rect 3472 -2632 3478 -2506
rect 3512 -2632 3518 -2506
rect 3278 -2650 3420 -2644
rect 3278 -2784 3350 -2650
rect 3472 -2686 3518 -2632
rect 3566 -2506 3710 -2494
rect 3566 -2632 3574 -2506
rect 3608 -2632 3710 -2506
rect 3758 -2512 3816 -2508
rect 3756 -2520 3822 -2512
rect 3756 -2572 3762 -2520
rect 3814 -2572 3822 -2520
rect 3756 -2578 3822 -2572
rect 3902 -2596 3908 -2474
rect 3942 -2596 3948 -2470
rect 3998 -2470 4044 -2458
rect 4092 -2466 4158 -2343
rect 3998 -2588 4004 -2470
rect 3902 -2608 3948 -2596
rect 3994 -2596 4004 -2588
rect 4038 -2596 4044 -2470
rect 3566 -2642 3710 -2632
rect 3568 -2644 3614 -2642
rect 3472 -2700 3580 -2686
rect 3472 -2756 3492 -2700
rect 3554 -2756 3580 -2700
rect 3472 -2776 3580 -2756
rect 3278 -2830 3342 -2784
rect 3098 -2866 3144 -2854
rect 3098 -2940 3104 -2866
rect 2923 -3138 2969 -3126
rect 2826 -3190 2874 -3138
rect 2634 -3230 2874 -3190
rect 1749 -3268 2028 -3262
rect 2091 -3268 2103 -3260
rect 14 -3303 1387 -3301
rect 1642 -3303 1761 -3268
rect 14 -3356 1510 -3303
rect 1580 -3311 1761 -3303
rect 2016 -3303 2103 -3268
rect 2358 -3268 2370 -3260
rect 2522 -3262 2640 -3260
rect 2522 -3264 2894 -3262
rect 2924 -3264 2968 -3138
rect 3092 -3142 3104 -2940
rect 3138 -3142 3144 -2866
rect 3092 -3260 3144 -3142
rect 3186 -2866 3244 -2854
rect 3186 -3142 3192 -2866
rect 3226 -3000 3244 -2866
rect 3274 -2838 3342 -2830
rect 3274 -2890 3284 -2838
rect 3336 -2890 3342 -2838
rect 3274 -2896 3342 -2890
rect 3370 -2818 3420 -2812
rect 3370 -2830 3422 -2818
rect 3370 -2900 3382 -2830
rect 3226 -3040 3232 -3000
rect 3226 -3048 3286 -3040
rect 3376 -3048 3382 -2900
rect 3278 -3100 3286 -3048
rect 3226 -3106 3286 -3100
rect 3352 -3056 3382 -3048
rect 3226 -3142 3232 -3106
rect 3352 -3108 3362 -3056
rect 3416 -3106 3422 -2830
rect 3414 -3108 3422 -3106
rect 3352 -3114 3422 -3108
rect 3376 -3118 3422 -3114
rect 3472 -2830 3518 -2776
rect 3472 -3106 3478 -2830
rect 3512 -3106 3518 -2830
rect 3472 -3118 3518 -3106
rect 3568 -2828 3614 -2818
rect 3568 -2830 3642 -2828
rect 3568 -3106 3574 -2830
rect 3608 -2836 3642 -2830
rect 3634 -2888 3642 -2836
rect 3608 -2894 3642 -2888
rect 3670 -2892 3710 -2642
rect 3994 -2698 4044 -2596
rect 4094 -2470 4140 -2466
rect 4094 -2596 4100 -2470
rect 4134 -2596 4140 -2470
rect 4094 -2608 4140 -2596
rect 4356 -2558 4408 -2341
rect 4356 -2684 4366 -2558
rect 4400 -2684 4408 -2558
rect 4356 -2696 4408 -2684
rect 4448 -2558 4494 -2546
rect 4448 -2684 4454 -2558
rect 4488 -2628 4494 -2558
rect 4488 -2684 4508 -2628
rect 4448 -2696 4508 -2684
rect 3994 -2718 4048 -2698
rect 3992 -2722 4280 -2718
rect 3992 -2724 4282 -2722
rect 3738 -2738 3812 -2726
rect 3738 -2790 3744 -2738
rect 3796 -2790 3812 -2738
rect 3992 -2730 4370 -2724
rect 3992 -2736 4376 -2730
rect 3992 -2772 4246 -2736
rect 3738 -2798 3812 -2790
rect 3994 -2804 4048 -2772
rect 4194 -2788 4246 -2772
rect 4298 -2752 4376 -2736
rect 4298 -2786 4330 -2752
rect 4364 -2786 4376 -2752
rect 4298 -2788 4376 -2786
rect 4194 -2804 4376 -2788
rect 3803 -2858 3849 -2846
rect 3608 -3106 3614 -2894
rect 3670 -3046 3718 -2892
rect 3568 -3118 3614 -3106
rect 3646 -3054 3718 -3046
rect 3646 -3106 3656 -3054
rect 3708 -3106 3718 -3054
rect 3646 -3112 3718 -3106
rect 3803 -3110 3809 -2858
rect 3186 -3154 3232 -3142
rect 3792 -3134 3809 -3110
rect 3843 -3110 3849 -2858
rect 3899 -2858 3945 -2846
rect 3994 -2856 4044 -2804
rect 3843 -3134 3850 -3110
rect 3332 -3164 3390 -3162
rect 3324 -3172 3394 -3164
rect 3324 -3224 3334 -3172
rect 3386 -3224 3394 -3172
rect 3792 -3180 3850 -3134
rect 3899 -3134 3905 -2858
rect 3939 -3134 3945 -2858
rect 3899 -3144 3945 -3134
rect 3995 -2858 4041 -2856
rect 3995 -3134 4001 -2858
rect 4035 -3134 4041 -2858
rect 3324 -3230 3394 -3224
rect 2522 -3268 2968 -3264
rect 3027 -3266 3306 -3260
rect 3027 -3268 3039 -3266
rect 2358 -3303 2627 -3268
rect 2016 -3311 2627 -3303
rect 2882 -3309 3039 -3268
rect 3294 -3268 3306 -3266
rect 3355 -3268 3634 -3262
rect 3794 -3268 3846 -3180
rect 3898 -3198 3946 -3144
rect 3995 -3146 4041 -3134
rect 4091 -2858 4137 -2846
rect 4091 -3134 4097 -2858
rect 4131 -3134 4137 -2858
rect 4091 -3146 4137 -3134
rect 4187 -2858 4233 -2846
rect 4187 -3134 4193 -2858
rect 4227 -3134 4233 -2858
rect 4456 -2862 4508 -2696
rect 4362 -2874 4408 -2862
rect 4362 -2948 4368 -2874
rect 4187 -3146 4233 -3134
rect 4090 -3198 4138 -3146
rect 3898 -3238 4138 -3198
rect 4188 -3268 4232 -3146
rect 4356 -3150 4368 -2948
rect 4402 -3150 4408 -2874
rect 4356 -3268 4408 -3150
rect 4450 -2874 4508 -2862
rect 4450 -3150 4456 -2874
rect 4490 -3008 4508 -2874
rect 4490 -3048 4496 -3008
rect 4490 -3056 4550 -3048
rect 4542 -3108 4550 -3056
rect 4490 -3114 4550 -3108
rect 4490 -3150 4496 -3114
rect 4450 -3162 4496 -3150
rect 4530 -3268 4652 -3258
rect 3294 -3309 3367 -3268
rect 2882 -3311 3367 -3309
rect 3622 -3274 4652 -3268
rect 3622 -3276 4303 -3274
rect 3622 -3311 3891 -3276
rect 1580 -3319 3891 -3311
rect 4146 -3317 4303 -3276
rect 4558 -3317 4652 -3274
rect 4146 -3319 4652 -3317
rect 1580 -3356 4652 -3319
rect 14 -3382 4652 -3356
rect 4530 -3408 4652 -3382
<< via1 >>
rect 1512 1032 1580 1088
rect 40 176 130 258
rect 2100 -62 2184 42
rect 66 -922 142 -856
rect 1510 -1146 1586 -1090
rect 40 -2020 132 -1922
rect 2094 -2278 2184 -2206
rect 2094 -2282 2104 -2278
rect 2104 -2282 2184 -2278
rect 626 -2558 678 -2492
rect 744 -2664 762 -2616
rect 762 -2664 796 -2616
rect 796 -2664 802 -2616
rect 744 -2668 802 -2664
rect 588 -2728 664 -2712
rect 588 -2762 604 -2728
rect 604 -2762 638 -2728
rect 638 -2762 664 -2728
rect 588 -2782 664 -2762
rect 2154 -2376 2206 -2368
rect 1536 -2618 1588 -2610
rect 1536 -2652 1546 -2618
rect 1546 -2652 1580 -2618
rect 1580 -2652 1588 -2618
rect 1536 -2662 1588 -2652
rect 2154 -2410 2162 -2376
rect 2162 -2410 2196 -2376
rect 2196 -2410 2206 -2376
rect 2154 -2420 2206 -2410
rect 948 -2798 1000 -2746
rect 1586 -2766 1638 -2714
rect 626 -3002 692 -2942
rect 1550 -2850 1602 -2838
rect 1550 -2884 1558 -2850
rect 1558 -2884 1592 -2850
rect 1592 -2884 1602 -2850
rect 1550 -2890 1602 -2884
rect 2496 -2518 2548 -2510
rect 2496 -2552 2506 -2518
rect 2506 -2552 2540 -2518
rect 2540 -2552 2548 -2518
rect 2496 -2562 2548 -2552
rect 2228 -2748 2290 -2692
rect 1712 -3176 1764 -3172
rect 1712 -3210 1720 -3176
rect 1720 -3210 1754 -3176
rect 1754 -3210 1764 -3176
rect 1712 -3224 1764 -3210
rect 2020 -2882 2072 -2830
rect 2098 -3098 2118 -3048
rect 2118 -3098 2150 -3048
rect 2098 -3100 2150 -3098
rect 2318 -2880 2344 -2828
rect 2344 -2880 2370 -2828
rect 3516 -2388 3568 -2380
rect 3516 -2422 3524 -2388
rect 3524 -2422 3558 -2388
rect 3558 -2422 3568 -2388
rect 3516 -2432 3568 -2422
rect 2480 -2740 2532 -2730
rect 2480 -2774 2494 -2740
rect 2494 -2774 2528 -2740
rect 2528 -2774 2532 -2740
rect 2480 -2782 2532 -2774
rect 2982 -2780 3034 -2728
rect 2392 -3098 2444 -3046
rect 2070 -3172 2122 -3164
rect 2070 -3206 2080 -3172
rect 2080 -3206 2114 -3172
rect 2114 -3206 2122 -3172
rect 2070 -3216 2122 -3206
rect 3762 -2526 3814 -2520
rect 3762 -2560 3770 -2526
rect 3770 -2560 3804 -2526
rect 3804 -2560 3814 -2526
rect 3762 -2572 3814 -2560
rect 3492 -2756 3554 -2700
rect 1510 -3303 1580 -3290
rect 1510 -3356 1580 -3303
rect 3284 -2890 3336 -2838
rect 3226 -3100 3278 -3048
rect 3362 -3106 3382 -3056
rect 3382 -3106 3414 -3056
rect 3362 -3108 3414 -3106
rect 3582 -2888 3608 -2836
rect 3608 -2888 3634 -2836
rect 3744 -2748 3796 -2738
rect 3744 -2782 3758 -2748
rect 3758 -2782 3792 -2748
rect 3792 -2782 3796 -2748
rect 3744 -2790 3796 -2782
rect 4246 -2788 4298 -2736
rect 3656 -3106 3708 -3054
rect 3334 -3180 3386 -3172
rect 3334 -3214 3344 -3180
rect 3344 -3214 3378 -3180
rect 3378 -3214 3386 -3180
rect 3334 -3224 3386 -3214
rect 4490 -3108 4542 -3056
<< metal2 >>
rect 1500 1088 1596 1098
rect 1500 1032 1512 1088
rect 1580 1032 1596 1088
rect 1500 1018 1596 1032
rect 3722 1008 3838 1020
rect 3722 938 3748 1008
rect 3812 938 3838 1008
rect 3722 918 3838 938
rect 12 258 154 264
rect 12 176 40 258
rect 130 176 154 258
rect 12 166 154 176
rect 2076 42 2216 58
rect 2076 -62 2100 42
rect 2184 -62 2216 42
rect 2076 -70 2216 -62
rect 44 -856 166 -840
rect 44 -922 66 -856
rect 142 -922 166 -856
rect 44 -938 166 -922
rect 3732 -944 3818 -928
rect 3732 -1002 3744 -944
rect 3802 -1002 3818 -944
rect 3732 -1018 3818 -1002
rect 1476 -1090 1632 -1082
rect 1476 -1146 1510 -1090
rect 1586 -1146 1632 -1090
rect 1476 -1162 1632 -1146
rect 3718 -1258 3804 -1242
rect 3718 -1316 3730 -1258
rect 3788 -1316 3804 -1258
rect 3718 -1332 3804 -1316
rect -2 -1598 122 -1588
rect -2 -1632 132 -1598
rect -2 -1706 36 -1632
rect 102 -1706 132 -1632
rect -2 -1740 132 -1706
rect 16 -1922 164 -1896
rect 16 -2020 40 -1922
rect 132 -2020 164 -1922
rect 2982 -1912 3056 -1900
rect 2982 -1970 2992 -1912
rect 3050 -1970 3056 -1912
rect 2982 -1986 3056 -1970
rect 16 -2048 164 -2020
rect 2060 -2206 2212 -2190
rect 2060 -2282 2094 -2206
rect 2184 -2282 2212 -2206
rect 2060 -2306 2212 -2282
rect 2020 -2362 2452 -2350
rect 3284 -2362 3716 -2358
rect 2020 -2368 3716 -2362
rect 2020 -2420 2154 -2368
rect 2206 -2380 3716 -2368
rect 2206 -2420 3516 -2380
rect 2020 -2422 3516 -2420
rect 2020 -2430 2452 -2422
rect 3284 -2432 3516 -2422
rect 3568 -2432 3716 -2380
rect 3284 -2438 3716 -2432
rect 14 -2444 152 -2440
rect 3496 -2442 3584 -2438
rect 14 -2480 678 -2444
rect 14 -2560 44 -2480
rect 114 -2492 686 -2480
rect 114 -2558 626 -2492
rect 678 -2558 686 -2492
rect 114 -2560 686 -2558
rect 14 -2566 686 -2560
rect 16 -2576 686 -2566
rect 1702 -2508 4622 -2492
rect 1702 -2510 2960 -2508
rect 1702 -2562 2496 -2510
rect 2548 -2562 2960 -2510
rect 1702 -2566 2960 -2562
rect 3018 -2520 4622 -2508
rect 3018 -2566 3762 -2520
rect 1702 -2572 3762 -2566
rect 3814 -2572 4622 -2520
rect 16 -2582 678 -2576
rect 1702 -2582 4622 -2572
rect 806 -2612 1536 -2610
rect 736 -2616 1536 -2612
rect 736 -2666 744 -2616
rect 738 -2668 744 -2666
rect 802 -2662 1536 -2616
rect 1588 -2662 1616 -2610
rect 802 -2666 1616 -2662
rect 802 -2668 808 -2666
rect 738 -2670 808 -2668
rect 1504 -2674 1616 -2666
rect 2416 -2680 2544 -2668
rect 2210 -2692 2544 -2680
rect 3680 -2688 3808 -2676
rect 582 -2712 680 -2704
rect 582 -2782 588 -2712
rect 664 -2782 680 -2712
rect 1580 -2714 1756 -2706
rect 582 -2792 680 -2782
rect 910 -2746 1048 -2728
rect 910 -2798 948 -2746
rect 1000 -2798 1048 -2746
rect 1580 -2766 1586 -2714
rect 1638 -2766 1756 -2714
rect 2210 -2748 2228 -2692
rect 2290 -2730 2544 -2692
rect 3474 -2700 3808 -2688
rect 3270 -2710 3342 -2708
rect 2290 -2748 2480 -2730
rect 2210 -2760 2480 -2748
rect 1580 -2778 1756 -2766
rect 910 -2816 1048 -2798
rect 1684 -2812 1754 -2778
rect 2416 -2782 2480 -2760
rect 2532 -2782 2544 -2730
rect 2416 -2790 2544 -2782
rect 2962 -2728 3342 -2710
rect 2962 -2780 2982 -2728
rect 3034 -2780 3342 -2728
rect 3474 -2756 3492 -2700
rect 3554 -2738 3808 -2700
rect 3554 -2756 3744 -2738
rect 3474 -2768 3744 -2756
rect 2962 -2802 3342 -2780
rect 3680 -2790 3744 -2768
rect 3796 -2790 3808 -2738
rect 3680 -2798 3808 -2790
rect 4226 -2736 4602 -2718
rect 4226 -2788 4246 -2736
rect 4298 -2788 4602 -2736
rect 1684 -2814 2078 -2812
rect 910 -2826 1628 -2816
rect 918 -2838 1628 -2826
rect 918 -2882 1550 -2838
rect 1542 -2890 1550 -2882
rect 1602 -2882 1628 -2838
rect 1684 -2828 2380 -2814
rect 1684 -2830 2318 -2828
rect 1684 -2882 2020 -2830
rect 2072 -2880 2318 -2830
rect 2370 -2880 2380 -2828
rect 2072 -2882 2380 -2880
rect 1602 -2890 1616 -2882
rect 1542 -2898 1616 -2890
rect 1684 -2892 2380 -2882
rect 3270 -2822 3342 -2802
rect 4226 -2810 4602 -2788
rect 3270 -2836 3644 -2822
rect 3270 -2838 3582 -2836
rect 3270 -2890 3284 -2838
rect 3336 -2888 3582 -2838
rect 3634 -2888 3644 -2836
rect 3336 -2890 3644 -2888
rect 1684 -2900 2078 -2892
rect 3270 -2900 3644 -2890
rect 4294 -2936 4358 -2810
rect 788 -2938 4358 -2936
rect 612 -2942 4358 -2938
rect 612 -3002 626 -2942
rect 692 -3000 4358 -2942
rect 692 -3002 4346 -3000
rect 612 -3008 836 -3002
rect 2384 -3038 3292 -3034
rect 2078 -3046 3292 -3038
rect 3648 -3046 4556 -3042
rect 2078 -3048 2392 -3046
rect 2078 -3100 2098 -3048
rect 2150 -3098 2392 -3048
rect 2444 -3048 3292 -3046
rect 2444 -3098 3226 -3048
rect 2150 -3100 3226 -3098
rect 3278 -3100 3292 -3048
rect 2078 -3110 3292 -3100
rect 2384 -3114 3292 -3110
rect 3342 -3054 4556 -3046
rect 3342 -3056 3656 -3054
rect 3342 -3108 3362 -3056
rect 3414 -3106 3656 -3056
rect 3708 -3056 4556 -3054
rect 3708 -3106 4490 -3056
rect 3414 -3108 4490 -3106
rect 4542 -3108 4556 -3056
rect 3342 -3118 4556 -3108
rect 3648 -3122 4556 -3118
rect 2040 -3154 2474 -3142
rect 3304 -3152 3738 -3150
rect 3304 -3154 4630 -3152
rect 2028 -3156 4630 -3154
rect 1696 -3164 4630 -3156
rect 1696 -3172 2070 -3164
rect 1696 -3224 1712 -3172
rect 1764 -3216 2070 -3172
rect 2122 -3172 4630 -3164
rect 2122 -3216 3334 -3172
rect 1764 -3224 3334 -3216
rect 3386 -3224 3736 -3172
rect 1696 -3230 3736 -3224
rect 3794 -3230 4630 -3172
rect 1696 -3234 4630 -3230
rect 1696 -3236 3810 -3234
rect 2028 -3240 3810 -3236
rect 3724 -3246 3810 -3240
rect 1490 -3290 1604 -3280
rect 1490 -3356 1510 -3290
rect 1580 -3356 1604 -3290
rect 1490 -3382 1604 -3356
<< via2 >>
rect 1512 1032 1580 1088
rect 3748 938 3812 1008
rect 40 176 130 258
rect 2986 252 3044 310
rect 2100 -62 2184 42
rect 2984 -334 3042 -276
rect 48 -604 108 -548
rect 68 -918 138 -860
rect 3744 -1002 3802 -944
rect 1510 -1146 1586 -1090
rect 3730 -1316 3788 -1258
rect 36 -1706 102 -1632
rect 40 -2020 132 -1922
rect 2992 -1970 3050 -1912
rect 2094 -2282 2184 -2206
rect 44 -2560 114 -2480
rect 2960 -2566 3018 -2508
rect 3736 -3230 3794 -3172
rect 1510 -3356 1580 -3290
<< metal3 >>
rect 1490 1088 1608 1118
rect 1490 1032 1512 1088
rect 1580 1070 1608 1088
rect 1580 1032 1612 1070
rect 1490 1030 1612 1032
rect 2 270 168 300
rect 2 258 170 270
rect 2 176 40 258
rect 130 176 170 258
rect 2 -548 170 176
rect 2 -604 48 -548
rect 108 -604 170 -548
rect 2 -614 170 -604
rect 74 -620 170 -614
rect 16 -848 156 -828
rect 14 -860 156 -848
rect 12 -918 68 -860
rect 138 -898 156 -860
rect 138 -918 154 -898
rect 12 -1632 154 -918
rect 12 -1706 36 -1632
rect 102 -1706 154 -1632
rect 12 -1720 154 -1706
rect 1492 -1090 1612 1030
rect 1492 -1146 1510 -1090
rect 1586 -1146 1612 -1090
rect 16 -1922 164 -1896
rect 16 -2020 40 -1922
rect 132 -2020 164 -1922
rect 16 -2048 164 -2020
rect 18 -2362 164 -2048
rect 18 -2480 172 -2362
rect 18 -2560 44 -2480
rect 114 -2560 172 -2480
rect 18 -2570 172 -2560
rect 18 -2580 164 -2570
rect -12 -3382 130 -3222
rect 1492 -3290 1612 -1146
rect 1492 -3356 1510 -3290
rect 1580 -3356 1612 -3290
rect 1492 -3388 1612 -3356
rect 2080 42 2200 1100
rect 3706 1008 3886 1020
rect 3706 938 3748 1008
rect 3812 938 3886 1008
rect 2080 -62 2100 42
rect 2184 -62 2200 42
rect 2080 -2206 2200 -62
rect 2946 310 3122 382
rect 2946 252 2986 310
rect 3044 252 3122 310
rect 2946 -276 3122 252
rect 2946 -334 2984 -276
rect 3042 -334 3122 -276
rect 2946 -378 3122 -334
rect 2080 -2282 2094 -2206
rect 2184 -2282 2200 -2206
rect 2944 -838 3122 -378
rect 3706 -436 3886 938
rect 2944 -1912 3078 -838
rect 2944 -1970 2992 -1912
rect 3050 -1970 3078 -1912
rect 2944 -2254 3078 -1970
rect 3700 -944 3892 -436
rect 3700 -1002 3744 -944
rect 3802 -1002 3892 -944
rect 3700 -1258 3892 -1002
rect 3700 -1316 3730 -1258
rect 3788 -1316 3892 -1258
rect 3700 -2254 3892 -1316
rect 2080 -3358 2200 -2282
rect 2922 -2508 3098 -2254
rect 2922 -2566 2960 -2508
rect 3018 -2566 3098 -2508
rect 2922 -3070 3098 -2566
rect 3682 -3070 3892 -2254
rect 3700 -3172 3892 -3070
rect 3700 -3230 3736 -3172
rect 3794 -3230 3892 -3172
rect 3700 -3378 3892 -3230
use bctr  bctr_0 cells
timestamp 1710564995
transform 1 0 1702 0 1 -2212
box -1704 -6 2946 1082
use bctr  bctr_2
timestamp 1710564995
transform 1 0 1694 0 1 12
box -1704 -6 2946 1082
use bctr  bctr_3
timestamp 1710564995
transform 1 0 1708 0 -1 -38
box -1704 -6 2946 1082
<< labels >>
rlabel space 1661 -93 2100 67 1 gnd
rlabel space 2532 1002 2650 1120 1 V
rlabel space 798 678 4356 744 1 Q1
rlabel space -10 516 324 590 1 CE
rlabel space 3396 892 3748 982 1 clk
rlabel space 812 -770 4370 -704 1 Q2
rlabel space 4264 -1746 4316 -1694 1 Q3
rlabel metal2 4298 -2810 4602 -2718 1 Q4
<< end >>
