magic
tech sky130A
magscale 1 2
timestamp 1709929695
<< nwell >>
rect 548 628 610 632
<< poly >>
rect 92 426 122 596
rect 188 426 218 598
rect 466 284 496 602
<< metal1 >>
rect 138 908 172 1002
rect 288 984 348 1034
rect 420 904 454 996
rect 548 628 610 632
rect 42 538 76 616
rect 234 538 268 616
rect 508 604 610 628
rect 42 506 474 538
rect 234 410 268 506
rect 582 464 610 604
rect 508 430 610 464
rect 508 266 542 430
rect 42 36 76 132
rect 280 6 354 50
rect 420 38 454 130
use grid  grid_0
timestamp 1678218586
transform 1 0 373 0 1 10
box -61 -10 259 1053
use grid  grid_1
timestamp 1678218586
transform 1 0 61 0 1 10
box -61 -10 259 1053
use sky130_fd_pr__nfet_01v8_NDWVGB  sky130_fd_pr__nfet_01v8_NDWVGB_0
timestamp 1709840560
transform 1 0 481 0 1 195
box -73 -101 73 101
use sky130_fd_pr__nfet_01v8_PLCS8W  sky130_fd_pr__nfet_01v8_PLCS8W_0
timestamp 1709840337
transform 1 0 155 0 1 262
box -125 -176 125 176
use sky130_fd_pr__pfet_01v8_52K3FE  sky130_fd_pr__pfet_01v8_52K3FE_0
timestamp 1709840560
transform 1 0 481 0 1 766
box -109 -212 109 212
use sky130_fd_pr__pfet_01v8_527QMA  sky130_fd_pr__pfet_01v8_527QMA_0
timestamp 1709840706
transform 1 0 155 0 1 760
box -161 -212 161 212
use via_m1_p  via_m1_p_0
timestamp 1646951168
transform 1 0 446 0 1 494
box 0 0 68 68
<< labels >>
rlabel metal1 280 6 354 50 1 vss
rlabel metal1 288 984 348 1034 1 vdd
rlabel space 92 412 122 610 1 a
rlabel space 188 412 218 610 1 b
rlabel metal1 508 430 610 464 1 out
<< end >>
