magic
tech sky130A
magscale 1 2
timestamp 1710542385
<< nwell >>
rect -1696 1052 -770 1076
rect -78 1074 290 1082
rect -78 1070 306 1074
rect -78 1068 304 1070
rect -1202 1048 -796 1052
rect -1202 1034 -798 1048
rect -1202 1016 -640 1034
rect -1202 990 -784 1016
rect -1202 776 -798 990
rect -1202 750 -980 776
rect -1202 660 -974 750
rect -896 732 -798 776
rect -14 732 304 1068
rect -896 728 304 732
rect -1202 652 -980 660
rect -896 652 -798 728
rect -1202 560 -798 652
rect -1202 534 -790 560
rect -14 556 304 728
rect -1202 484 -1120 534
rect -1080 474 -790 534
rect -16 520 994 556
rect -16 519 274 520
rect -20 514 274 519
rect -22 508 274 514
rect 420 508 994 520
rect -22 496 218 508
rect -22 490 280 496
rect 512 490 994 508
rect 512 482 698 490
<< poly >>
rect -1052 482 -888 494
rect -1052 460 -838 482
rect -916 456 -838 460
<< metal1 >>
rect -1008 1024 -640 1034
rect -1030 1016 -640 1024
rect -1030 994 -946 1016
rect -1072 750 -1002 856
rect -1072 732 -974 750
rect -1072 672 -1058 732
rect -992 672 -974 732
rect -1072 660 -974 672
rect -1072 440 -1002 660
rect -1064 296 -1002 306
rect -1064 164 -990 296
rect -1064 102 -858 164
rect -1014 4 -621 52
rect -47 4 135 55
<< via1 >>
rect -1058 672 -992 732
<< metal2 >>
rect -1636 880 44 952
rect -1072 732 -848 738
rect -1072 672 -1058 732
rect -992 730 2662 732
rect -992 672 2674 730
rect -1072 668 2674 672
rect -896 666 2674 668
rect -1704 504 -1372 578
rect 0 508 70 624
rect -104 436 72 508
rect 2610 448 2674 666
rect 12 310 50 312
rect 10 294 50 310
rect -1666 292 50 294
rect -1666 244 52 292
rect -1656 230 52 244
rect -1656 220 50 230
rect -1656 218 18 220
use and  and_0 cells
timestamp 1710542385
transform -1 0 -1066 0 1 -6
box -62 0 632 1063
use ffdr3  ffdr3_0 cells
timestamp 1710538400
transform 1 0 322 0 1 2
box -322 -2 2624 1079
use xor  xor_0 xor
timestamp 1710539684
transform 1 0 -662 0 1 0
box -386 -4 652 1074
<< end >>
