magic
tech sky130A
magscale 1 2
timestamp 1710257160
<< nwell >>
rect -708 1135 336 1136
rect -708 1134 944 1135
rect -708 1126 1688 1134
rect -426 602 86 1126
rect -426 588 -340 602
rect -436 586 -340 588
rect -284 588 86 602
rect -284 586 276 588
rect -436 582 276 586
rect -436 552 -264 582
rect -240 554 -116 582
rect -30 550 276 582
rect 316 558 1688 1126
rect 916 550 1688 558
rect 1322 548 1628 550
<< nmos >>
rect 766 332 796 482
rect 458 176 488 326
rect 1116 234 1146 384
rect 1212 234 1242 384
rect 1510 168 1540 318
<< pmos >>
rect 458 686 488 986
rect 768 648 798 948
rect 1017 622 1047 922
rect 1113 622 1143 922
rect 1209 622 1239 922
rect 1305 622 1335 922
rect 1510 678 1540 978
<< ndiff >>
rect 708 470 766 482
rect 708 344 720 470
rect 754 344 766 470
rect 708 332 766 344
rect 796 470 854 482
rect 796 344 808 470
rect 842 344 854 470
rect 796 332 854 344
rect 400 314 458 326
rect 400 188 412 314
rect 446 188 458 314
rect 400 176 458 188
rect 488 314 546 326
rect 488 188 500 314
rect 534 188 546 314
rect 1054 372 1116 384
rect 1054 246 1066 372
rect 1100 246 1116 372
rect 1054 234 1116 246
rect 1146 372 1212 384
rect 1146 246 1162 372
rect 1196 246 1212 372
rect 1146 234 1212 246
rect 1242 372 1304 384
rect 1242 246 1258 372
rect 1292 246 1304 372
rect 1242 234 1304 246
rect 1452 306 1510 318
rect 488 176 546 188
rect 1452 180 1464 306
rect 1498 180 1510 306
rect 1452 168 1510 180
rect 1540 306 1598 318
rect 1540 180 1552 306
rect 1586 180 1598 306
rect 1540 168 1598 180
<< pdiff >>
rect 400 974 458 986
rect 400 698 412 974
rect 446 698 458 974
rect 400 686 458 698
rect 488 974 546 986
rect 488 698 500 974
rect 534 698 546 974
rect 488 686 546 698
rect 710 936 768 948
rect 710 660 722 936
rect 756 660 768 936
rect 710 648 768 660
rect 798 936 856 948
rect 798 660 810 936
rect 844 660 856 936
rect 1452 966 1510 978
rect 798 648 856 660
rect 955 910 1017 922
rect 955 634 967 910
rect 1001 634 1017 910
rect 955 622 1017 634
rect 1047 910 1113 922
rect 1047 634 1063 910
rect 1097 634 1113 910
rect 1047 622 1113 634
rect 1143 910 1209 922
rect 1143 634 1159 910
rect 1193 634 1209 910
rect 1143 622 1209 634
rect 1239 910 1305 922
rect 1239 634 1255 910
rect 1289 634 1305 910
rect 1239 622 1305 634
rect 1335 910 1397 922
rect 1335 634 1351 910
rect 1385 634 1397 910
rect 1452 690 1464 966
rect 1498 690 1510 966
rect 1452 678 1510 690
rect 1540 966 1598 978
rect 1540 690 1552 966
rect 1586 690 1598 966
rect 1540 678 1598 690
rect 1335 622 1397 634
<< ndiffc >>
rect 720 344 754 470
rect 808 344 842 470
rect 412 188 446 314
rect 500 188 534 314
rect 1066 246 1100 372
rect 1162 246 1196 372
rect 1258 246 1292 372
rect 1464 180 1498 306
rect 1552 180 1586 306
<< pdiffc >>
rect 412 698 446 974
rect 500 698 534 974
rect 722 660 756 936
rect 810 660 844 936
rect 967 634 1001 910
rect 1063 634 1097 910
rect 1159 634 1193 910
rect 1255 634 1289 910
rect 1351 634 1385 910
rect 1464 690 1498 966
rect 1552 690 1586 966
<< psubdiff >>
rect 357 82 381 116
rect 581 82 605 116
rect 661 82 685 116
rect 885 82 909 116
rect 1053 74 1077 108
rect 1277 74 1301 108
rect 1405 74 1429 108
rect 1629 74 1653 108
<< nsubdiff >>
rect 366 1098 614 1099
rect 366 1064 415 1098
rect 562 1064 614 1098
rect 366 1063 614 1064
rect 684 1098 932 1099
rect 684 1064 733 1098
rect 880 1064 932 1098
rect 684 1063 932 1064
rect 1052 1090 1300 1091
rect 1052 1056 1101 1090
rect 1248 1056 1300 1090
rect 1052 1055 1300 1056
rect 1404 1090 1652 1091
rect 1404 1056 1453 1090
rect 1600 1056 1652 1090
rect 1404 1055 1652 1056
<< psubdiffcont >>
rect 381 82 581 116
rect 685 82 885 116
rect 1077 74 1277 108
rect 1429 74 1629 108
<< nsubdiffcont >>
rect 415 1064 562 1098
rect 733 1064 880 1098
rect 1101 1056 1248 1090
rect 1453 1056 1600 1090
<< poly >>
rect -336 998 -20 1026
rect -336 996 -16 998
rect -336 950 -304 996
rect -52 942 -16 996
rect 458 986 488 1012
rect 1016 996 1332 1024
rect 1016 994 1336 996
rect 768 948 798 974
rect 1016 948 1048 994
rect 458 660 488 686
rect 1017 922 1047 948
rect 1113 922 1143 952
rect 1209 922 1239 948
rect 1300 940 1336 994
rect 1510 978 1540 1004
rect 1305 922 1335 940
rect 768 630 798 648
rect -846 598 -568 604
rect 766 602 798 630
rect 1510 652 1540 678
rect -848 572 -566 598
rect -342 556 -300 600
rect -144 598 -112 600
rect -450 498 -300 556
rect -240 554 -112 598
rect -238 438 -200 554
rect -48 518 -16 598
rect 506 596 798 602
rect 1017 598 1047 622
rect 504 570 798 596
rect -48 442 -10 518
rect 766 504 798 570
rect 1010 554 1052 598
rect 1113 596 1143 622
rect 1209 598 1239 622
rect 1208 596 1240 598
rect 1305 596 1335 622
rect 766 482 796 504
rect 902 496 1052 554
rect 1112 552 1240 596
rect -366 410 -200 438
rect -140 412 -10 442
rect -366 408 -230 410
rect -366 398 -326 408
rect -442 284 -326 398
rect 458 326 488 352
rect 1114 436 1152 552
rect 1304 516 1336 596
rect 1304 440 1342 516
rect 986 408 1152 436
rect 1212 410 1342 440
rect 986 406 1146 408
rect 986 396 1026 406
rect 766 306 796 332
rect 910 282 1026 396
rect 1116 384 1146 406
rect 1212 384 1242 410
rect 1510 318 1540 344
rect 1116 208 1146 234
rect 1212 208 1242 234
rect 458 150 488 176
rect 1510 142 1540 168
<< locali >>
rect 357 1103 623 1106
rect 357 1060 363 1103
rect 618 1060 623 1103
rect 357 1056 623 1060
rect 675 1103 941 1106
rect 675 1060 681 1103
rect 936 1060 941 1103
rect 675 1056 941 1060
rect 1043 1095 1309 1098
rect 1043 1052 1049 1095
rect 1304 1052 1309 1095
rect 1043 1048 1309 1052
rect 1395 1095 1661 1098
rect 1395 1052 1401 1095
rect 1656 1052 1661 1095
rect 1395 1048 1661 1052
rect 412 974 446 990
rect 412 682 446 698
rect 500 974 534 990
rect 1464 966 1498 982
rect 500 682 534 698
rect 722 936 756 952
rect 722 644 756 660
rect 810 936 844 952
rect 810 644 844 660
rect 967 910 1001 926
rect 967 618 1001 634
rect 1063 910 1097 926
rect 1063 618 1097 634
rect 1159 910 1193 926
rect 1159 618 1193 634
rect 1255 910 1289 926
rect 1255 618 1289 634
rect 1351 910 1385 926
rect 1464 674 1498 690
rect 1552 966 1586 982
rect 1552 674 1586 690
rect 1351 618 1385 634
rect 720 470 754 486
rect 412 314 446 330
rect 412 172 446 188
rect 500 314 534 330
rect 720 328 754 344
rect 808 470 842 486
rect 808 328 842 344
rect 1066 372 1100 388
rect 1066 230 1100 246
rect 1162 372 1196 388
rect 1162 230 1196 246
rect 1258 372 1292 388
rect 1258 230 1292 246
rect 1464 306 1498 322
rect 500 172 534 188
rect 1464 164 1498 180
rect 1552 306 1586 322
rect 1552 164 1586 180
<< viali >>
rect 363 1098 618 1103
rect 363 1064 415 1098
rect 415 1064 562 1098
rect 562 1064 618 1098
rect 363 1060 618 1064
rect 681 1098 936 1103
rect 681 1064 733 1098
rect 733 1064 880 1098
rect 880 1064 936 1098
rect 681 1060 936 1064
rect 1049 1090 1304 1095
rect 1049 1056 1101 1090
rect 1101 1056 1248 1090
rect 1248 1056 1304 1090
rect 1049 1052 1304 1056
rect 1401 1090 1656 1095
rect 1401 1056 1453 1090
rect 1453 1056 1600 1090
rect 1600 1056 1656 1090
rect 1401 1052 1656 1056
rect 412 698 446 974
rect 500 698 534 974
rect 722 660 756 936
rect 810 660 844 936
rect 967 634 1001 910
rect 1063 634 1097 910
rect 1159 634 1193 910
rect 1255 634 1289 910
rect 1351 634 1385 910
rect 1464 690 1498 966
rect 1552 690 1586 966
rect 720 344 754 470
rect 412 188 446 314
rect 808 344 842 470
rect 500 188 534 314
rect 1066 246 1100 372
rect 1162 246 1196 372
rect 1258 246 1292 372
rect 1464 180 1498 306
rect 1552 180 1586 306
rect 354 116 609 121
rect 354 82 381 116
rect 381 82 581 116
rect 581 82 609 116
rect 354 78 609 82
rect 658 116 913 121
rect 658 82 685 116
rect 685 82 885 116
rect 885 82 913 116
rect 658 78 913 82
rect 1050 108 1305 113
rect 1050 74 1077 108
rect 1077 74 1277 108
rect 1277 74 1305 108
rect 1050 70 1305 74
rect 1402 108 1657 113
rect 1402 74 1429 108
rect 1429 74 1629 108
rect 1629 74 1657 108
rect 1402 70 1657 74
<< metal1 >>
rect 328 1132 362 1134
rect 286 1126 410 1132
rect -992 1124 410 1126
rect -992 1120 1692 1124
rect -1018 1103 1692 1120
rect -1018 1060 363 1103
rect 618 1060 681 1103
rect 936 1095 1692 1103
rect 936 1060 1049 1095
rect -1018 1058 1049 1060
rect -1018 1046 -290 1058
rect -42 1050 38 1058
rect -1018 1040 -348 1046
rect -400 958 -348 1040
rect -296 976 -56 1016
rect -402 888 -344 958
rect -296 922 -248 976
rect -104 924 -56 976
rect -6 874 38 1050
rect 286 1052 1049 1058
rect 1304 1052 1401 1095
rect 1656 1056 1692 1095
rect 1656 1052 1668 1056
rect 286 1048 1668 1052
rect 286 1046 1316 1048
rect 1346 1046 1668 1048
rect 286 1044 1062 1046
rect 286 1038 1004 1044
rect 286 1036 410 1038
rect 406 974 452 986
rect 406 698 412 974
rect 446 698 452 974
rect 406 686 452 698
rect 494 974 540 986
rect 494 698 500 974
rect 534 698 540 974
rect 710 936 762 1038
rect 952 956 1004 1038
rect 1056 974 1296 1014
rect 710 734 722 936
rect 494 686 540 698
rect -200 582 -150 634
rect -1038 516 -912 574
rect -540 570 -380 576
rect -540 518 -444 570
rect -386 518 -380 570
rect -200 550 -146 582
rect 284 578 376 590
rect -540 510 -380 518
rect -202 546 86 550
rect -540 508 -388 510
rect -202 496 142 546
rect -200 476 -146 496
rect 76 494 142 496
rect 284 526 308 578
rect 366 572 376 578
rect 414 572 446 686
rect 366 526 446 572
rect 284 514 446 526
rect 284 490 376 514
rect -200 366 -150 476
rect -444 348 -374 352
rect -446 346 -374 348
rect -446 294 -438 346
rect -380 294 -374 346
rect 414 326 446 514
rect 500 326 532 686
rect 716 660 722 734
rect 756 660 762 936
rect 716 648 762 660
rect 804 936 850 948
rect 804 660 810 936
rect 844 794 850 936
rect 950 910 1008 956
rect 1056 920 1104 974
rect 1248 922 1296 974
rect 1346 922 1390 1046
rect 1458 966 1504 978
rect 950 886 967 910
rect 844 660 862 794
rect 804 648 862 660
rect 810 574 862 648
rect 961 634 967 886
rect 1001 886 1008 910
rect 1057 910 1103 920
rect 1001 634 1007 886
rect 961 622 1007 634
rect 1057 634 1063 910
rect 1097 634 1103 910
rect 1057 622 1103 634
rect 1153 910 1199 922
rect 1153 634 1159 910
rect 1193 634 1199 910
rect 1153 632 1199 634
rect 1249 910 1295 922
rect 1249 634 1255 910
rect 1289 634 1295 910
rect 1152 580 1202 632
rect 1249 622 1295 634
rect 1345 910 1391 922
rect 1345 634 1351 910
rect 1385 634 1391 910
rect 1458 690 1464 966
rect 1498 690 1504 966
rect 1458 678 1504 690
rect 1546 966 1592 978
rect 1546 690 1552 966
rect 1586 690 1592 966
rect 1546 678 1592 690
rect 1345 622 1391 634
rect 810 568 972 574
rect 810 516 908 568
rect 966 516 972 568
rect 1152 548 1206 580
rect 810 508 972 516
rect 1150 544 1438 548
rect 1466 544 1498 678
rect 810 506 964 508
rect 810 482 862 506
rect 1150 494 1498 544
rect 710 470 762 482
rect 710 344 720 470
rect 754 344 762 470
rect -446 288 -374 294
rect -444 286 -374 288
rect 406 314 452 326
rect -856 234 -704 242
rect -856 182 -772 234
rect -714 182 -704 234
rect -856 162 -704 182
rect -310 148 -252 252
rect -344 134 -252 148
rect -102 134 -36 244
rect 270 234 340 238
rect 202 232 340 234
rect 202 180 276 232
rect 334 180 340 232
rect 202 174 340 180
rect 406 188 412 314
rect 446 188 452 314
rect 406 176 452 188
rect 494 314 540 326
rect 494 188 500 314
rect 534 240 540 314
rect 534 232 650 240
rect 534 188 580 232
rect 494 180 580 188
rect 638 180 650 232
rect 494 176 650 180
rect 270 172 340 174
rect 498 164 650 176
rect 286 134 368 138
rect -1014 132 368 134
rect 710 132 762 344
rect 802 470 862 482
rect 802 344 808 470
rect 842 414 862 470
rect 1152 474 1206 494
rect 1428 492 1498 494
rect 842 344 848 414
rect 1060 372 1106 384
rect 908 346 978 350
rect 802 332 848 344
rect 906 344 978 346
rect 906 292 914 344
rect 972 292 978 344
rect 906 286 978 292
rect 908 284 978 286
rect 1060 250 1066 372
rect 1042 246 1066 250
rect 1100 246 1106 372
rect 1152 372 1202 474
rect 1152 364 1162 372
rect 1042 234 1106 246
rect 1156 246 1162 364
rect 1196 246 1202 372
rect 1156 234 1202 246
rect 1252 372 1298 384
rect 1252 246 1258 372
rect 1292 246 1298 372
rect 1466 318 1498 492
rect 1552 318 1584 678
rect 1252 242 1298 246
rect 1458 306 1504 318
rect 1042 146 1100 234
rect 1008 132 1100 146
rect 1250 132 1316 242
rect 1458 180 1464 306
rect 1498 180 1504 306
rect 1458 168 1504 180
rect 1546 306 1592 318
rect 1546 180 1552 306
rect 1586 232 1592 306
rect 1622 232 1692 236
rect 1586 230 1692 232
rect 1586 180 1628 230
rect 1546 178 1628 180
rect 1686 178 1692 230
rect 1546 172 1692 178
rect 1546 168 1592 172
rect 1622 170 1692 172
rect -1014 130 1666 132
rect -1022 121 1666 130
rect -1022 78 354 121
rect 609 78 658 121
rect 913 119 1666 121
rect 913 113 1669 119
rect 913 78 1050 113
rect -1022 70 1050 78
rect 1305 70 1402 113
rect 1657 70 1669 113
rect -1022 64 1669 70
rect -1022 60 1666 64
rect -688 58 -191 60
rect -376 56 -191 58
rect -160 56 7 60
rect 286 58 1666 60
rect 664 56 1161 58
rect 976 54 1161 56
rect 1192 54 1359 58
<< via1 >>
rect -444 518 -386 570
rect 308 526 366 578
rect -438 294 -380 346
rect 908 516 966 568
rect -772 182 -714 234
rect 276 180 334 232
rect 580 180 638 232
rect 914 292 972 344
rect 1628 178 1686 230
<< metal2 >>
rect 284 584 376 590
rect -460 578 376 584
rect -460 570 308 578
rect -460 518 -444 570
rect -386 526 308 570
rect 366 526 376 578
rect -386 518 376 526
rect -460 498 376 518
rect 284 490 376 498
rect 892 568 1684 582
rect 892 516 908 568
rect 966 516 1684 568
rect 892 496 1684 516
rect -508 360 328 362
rect -1036 358 328 360
rect 844 358 1680 360
rect -1036 346 1680 358
rect -1036 294 -438 346
rect -380 344 1680 346
rect -380 294 914 344
rect -1036 292 914 294
rect 972 292 1680 344
rect -1036 274 1680 292
rect 316 272 1680 274
rect -782 234 346 242
rect -782 182 -772 234
rect -714 232 346 234
rect -714 182 276 232
rect -782 180 276 182
rect 334 180 346 232
rect -782 170 346 180
rect 268 168 346 170
rect 570 232 1698 240
rect 570 180 580 232
rect 638 230 1698 232
rect 638 180 1628 230
rect 570 178 1628 180
rect 1686 178 1698 230
rect 570 168 1698 178
rect 1620 166 1698 168
use grid#0  grid_0 /foss/designs/EAMTA2024/EAMTA/mag/ffdr/nor
timestamp 1678218586
transform 1 0 -275 0 1 76
box -61 -10 259 1053
use inv  inv_0 /foss/designs/EAMTA2024/EAMTA/mag
timestamp 1710256097
transform 1 0 -728 0 1 74
box 0 0 320 1063
use passGate  passGate_0 /foss/designs/EAMTA2024/EAMTA/mag/passGate
timestamp 1710256097
transform 1 0 86 0 1 -190
box -70 256 250 1319
use passGate  passGate_1
timestamp 1710256097
transform 1 0 -966 0 1 -182
box -70 256 250 1319
use sky130_fd_pr__nfet_01v8_XUMWGH  sky130_fd_pr__nfet_01v8_XUMWGH_0 /foss/designs/EAMTA2024/EAMTA/mag/ffdr/nor
timestamp 1710120945
transform 1 0 -173 0 1 311
box -125 -101 125 101
use sky130_fd_pr__pfet_01v8_52FGJA  sky130_fd_pr__pfet_01v8_52FGJA_0
timestamp 1710120945
transform 1 0 -176 0 1 774
box -260 -192 262 202
use via_m1_p  via_m1_p_0 /foss/designs/EAMTA2024/EAMTA/mag
timestamp 1646951168
transform 1 0 486 0 1 548
box 0 0 68 68
use via_m1_p  via_m1_p_1
timestamp 1646951168
transform 1 0 898 0 1 506
box 0 0 68 68
use via_m1_p  via_m1_p_2
timestamp 1646951168
transform 1 0 910 0 1 284
box 0 0 68 68
use via_m1_p  via_m1_p_3
timestamp 1646951168
transform 1 0 -866 0 1 550
box 0 0 68 68
use via_m1_p  via_m1_p_4
timestamp 1646951168
transform 1 0 -454 0 1 508
box 0 0 68 68
use via_m1_p  via_m1_p_5
timestamp 1646951168
transform 1 0 -442 0 1 286
box 0 0 68 68
<< labels >>
rlabel space -646 552 58 1129 1 V
rlabel space -623 56 57 115 1 gnd
rlabel poly -424 304 -390 338 1 B
rlabel metal1 -202 496 86 550 1 out
rlabel via1 -436 526 -402 560 1 A
rlabel pmos 1510 834 1540 902 1 clk_1
rlabel nmos 1510 216 1540 267 1 clk_2
rlabel metal1 1552 294 1584 536 1 out
rlabel metal1 1466 294 1498 536 1 in
rlabel pmos 458 842 488 910 1 clk_1
rlabel nmos 458 224 488 275 1 clk_2
rlabel metal1 500 302 532 544 1 out
rlabel metal1 414 302 446 544 1 in
rlabel poly 766 504 798 630 1 in
rlabel metal1 710 102 762 482 1 gnd
rlabel nwell 710 734 762 1114 1 V
rlabel metal1 810 414 862 794 1 out
rlabel via1 916 524 950 558 1 A
rlabel metal1 1150 494 1438 548 1 out
rlabel poly 928 302 962 336 1 B
rlabel space 729 54 1409 113 1 gnd
rlabel space 706 550 1410 1127 1 V
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
