magic
tech sky130A
magscale 1 2
timestamp 1710560808
<< error_s >>
rect 94 534 124 574
rect 320 518 332 764
rect 320 510 574 518
<< nwell >>
rect -284 1068 596 1074
rect -284 1052 652 1068
rect -284 1032 18 1052
rect -284 982 22 1032
rect -284 970 18 982
rect 192 970 222 1052
rect 314 1040 652 1052
rect -284 930 222 970
rect -284 542 18 930
rect 92 886 124 930
rect 180 908 222 930
rect 186 888 222 908
rect 224 968 652 1040
rect 224 964 242 968
rect 280 964 652 968
rect 224 898 652 964
rect 260 896 652 898
rect 260 894 276 896
rect -284 530 -120 542
rect -116 530 18 542
rect -284 482 18 530
rect 94 502 124 532
rect 192 502 222 888
rect 286 886 316 896
rect 414 894 652 896
rect 462 510 652 894
rect 288 486 652 510
<< poly >>
rect 286 972 556 974
rect -224 964 218 966
rect -224 958 222 964
rect -348 944 222 958
rect -358 934 222 944
rect -358 918 -170 934
rect -358 786 -304 918
rect -224 910 -170 918
rect -218 874 -174 910
rect 180 908 222 934
rect 186 904 222 908
rect 286 944 594 972
rect 186 888 220 904
rect 286 896 324 944
rect 470 934 594 944
rect 286 886 316 896
rect 522 608 594 934
rect -216 500 -174 538
rect -304 464 -174 500
rect -216 424 -174 464
rect -120 488 -74 534
rect 94 488 124 532
rect -120 440 124 488
rect -116 424 124 440
rect -116 422 118 424
rect 190 412 220 556
rect 286 412 316 572
rect 382 476 412 570
rect 380 434 568 476
rect 380 418 586 434
rect 382 410 412 418
rect 502 342 586 418
rect -116 202 -82 230
rect -122 168 -82 202
rect -288 104 -82 168
rect -122 102 -82 104
<< metal1 >>
rect 14 1026 22 1032
rect -284 992 22 1026
rect 300 1022 470 1036
rect -164 852 -124 992
rect 14 982 22 992
rect -72 886 -30 944
rect -72 848 -28 886
rect 134 858 180 1004
rect 298 982 470 1022
rect 230 922 466 950
rect 230 854 276 922
rect 414 896 466 922
rect 414 894 468 896
rect 422 860 468 894
rect -72 846 -30 848
rect -282 398 -216 590
rect -78 538 -20 596
rect -96 528 2 538
rect -96 476 -74 528
rect -22 476 2 528
rect 38 532 84 560
rect 230 532 276 560
rect 38 504 276 532
rect 326 506 372 560
rect -96 452 2 476
rect 326 496 652 506
rect 326 472 564 496
rect -282 346 -278 398
rect -220 346 -216 398
rect -282 340 -216 346
rect -282 288 -230 340
rect -222 288 -216 340
rect -282 220 -216 288
rect -166 50 -114 258
rect -78 228 -20 452
rect 232 444 564 472
rect 616 444 652 496
rect 232 434 652 444
rect 232 404 274 434
rect 232 370 276 404
rect 14 50 22 52
rect 38 50 80 100
rect 424 54 464 100
rect -166 20 80 50
rect 296 48 464 54
rect -166 12 44 20
rect -166 6 -114 12
rect 14 0 22 12
rect 296 2 470 48
rect 420 -2 470 2
<< via1 >>
rect 528 568 580 620
rect -74 476 -22 528
rect -278 346 -220 398
rect 564 444 616 496
rect 514 340 566 392
<< metal2 >>
rect 520 620 594 628
rect 520 612 528 620
rect -104 568 528 612
rect 580 612 594 620
rect 580 568 606 612
rect -104 556 606 568
rect -112 546 606 556
rect -112 528 26 546
rect -112 476 -74 528
rect -22 476 26 528
rect -112 458 26 476
rect 558 496 628 502
rect 558 444 564 496
rect 616 444 628 496
rect 558 442 628 444
rect -284 398 -214 400
rect -284 396 -278 398
rect -286 346 -278 396
rect -220 396 -214 398
rect 482 396 594 404
rect -220 392 594 396
rect -220 346 514 392
rect -286 342 514 346
rect -216 340 514 342
rect 566 340 594 392
use grid#3  grid#3_0
timestamp 1709738583
transform 1 0 -261 0 1 6
box -61 -10 259 1053
use grid#3  grid_0
timestamp 1709738583
transform 1 0 61 0 1 10
box -61 -10 259 1053
use grid#3  grid_1
timestamp 1709738583
transform 1 0 393 0 1 12
box -61 -10 259 1053
use sky130_fd_pr__nfet_01v8_ND3UG5  sky130_fd_pr__nfet_01v8_ND3UG5_0
timestamp 1709927624
transform 1 0 253 0 1 250
box -221 -176 221 176
use sky130_fd_pr__nfet_01v8_XUMWGH  sky130_fd_pr__nfet_01v8_XUMWGH_0
timestamp 1710263695
transform 1 0 -147 0 1 331
box -125 -101 125 101
use sky130_fd_pr__pfet_01v8_52FGJA  sky130_fd_pr__pfet_01v8_52FGJA_0
timestamp 1710120945
transform 1 0 253 0 1 710
box -260 -192 262 202
use sky130_fd_pr__pfet_01v8_527QMA#1  sky130_fd_pr__pfet_01v8_527QMA_0
timestamp 1710106043
transform 1 0 -148 0 1 708
box -162 -186 162 186
use via_m1_p#2  via_m1_p_0
timestamp 1646951168
transform 1 0 -266 0 1 102
box 0 0 68 68
use via_m1_p#2  via_m1_p_1
timestamp 1646951168
transform 1 0 -386 0 1 798
box 0 0 68 68
use via_m1_p#2  via_m1_p_2
timestamp 1646951168
transform 1 0 506 0 1 330
box 0 0 68 68
use via_m1_p#2  via_m1_p_3
timestamp 1646951168
transform 1 0 518 0 1 562
box 0 0 68 68
<< labels >>
rlabel metal1 232 370 274 472 1 out
rlabel space 33 988 288 1031 1 V
rlabel nwell -246 922 -212 956 1 A
rlabel poly -248 120 -214 154 1 B
rlabel space 61 10 261 44 1 gnd
rlabel via1 524 348 558 382 1 nA
rlabel via1 528 568 580 620 1 nB
<< end >>
