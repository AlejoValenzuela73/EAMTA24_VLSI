magic
tech sky130A
magscale 1 2
timestamp 1710359923
<< nwell >>
rect 1852 1078 2172 1079
rect 1762 1077 2274 1078
rect 1762 1076 2584 1077
rect -44 1068 2584 1076
rect -48 488 1016 1068
rect 1216 500 2584 1068
rect 1216 496 2280 500
rect 1308 494 1648 496
rect 1308 490 1628 494
<< nmos >>
rect 1426 222 1456 372
rect 1522 222 1552 372
rect 1952 186 1982 336
rect 2048 186 2078 336
rect 2406 274 2436 424
<< pmos >>
rect 1426 546 1456 846
rect 1522 546 1552 846
rect 1853 574 1883 874
rect 1949 574 1979 874
rect 2045 574 2075 874
rect 2141 574 2171 874
rect 2408 590 2438 890
<< ndiff >>
rect 1364 360 1426 372
rect 1364 234 1376 360
rect 1410 234 1426 360
rect 1364 222 1426 234
rect 1456 360 1522 372
rect 1456 234 1472 360
rect 1506 234 1522 360
rect 1456 222 1522 234
rect 1552 360 1614 372
rect 1552 234 1568 360
rect 1602 234 1614 360
rect 2348 412 2406 424
rect 1890 324 1952 336
rect 1552 222 1614 234
rect 1890 198 1902 324
rect 1936 198 1952 324
rect 1890 186 1952 198
rect 1982 324 2048 336
rect 1982 198 1998 324
rect 2032 198 2048 324
rect 1982 186 2048 198
rect 2078 324 2140 336
rect 2078 198 2094 324
rect 2128 198 2140 324
rect 2348 286 2360 412
rect 2394 286 2406 412
rect 2348 274 2406 286
rect 2436 412 2494 424
rect 2436 286 2448 412
rect 2482 286 2494 412
rect 2436 274 2494 286
rect 2078 186 2140 198
<< pdiff >>
rect 2350 878 2408 890
rect 1791 862 1853 874
rect 1364 834 1426 846
rect 1364 558 1376 834
rect 1410 558 1426 834
rect 1364 546 1426 558
rect 1456 834 1522 846
rect 1456 558 1472 834
rect 1506 558 1522 834
rect 1456 546 1522 558
rect 1552 834 1614 846
rect 1552 558 1568 834
rect 1602 558 1614 834
rect 1791 586 1803 862
rect 1837 586 1853 862
rect 1791 574 1853 586
rect 1883 862 1949 874
rect 1883 586 1899 862
rect 1933 586 1949 862
rect 1883 574 1949 586
rect 1979 862 2045 874
rect 1979 586 1995 862
rect 2029 586 2045 862
rect 1979 574 2045 586
rect 2075 862 2141 874
rect 2075 586 2091 862
rect 2125 586 2141 862
rect 2075 574 2141 586
rect 2171 862 2233 874
rect 2171 586 2187 862
rect 2221 586 2233 862
rect 2350 602 2362 878
rect 2396 602 2408 878
rect 2350 590 2408 602
rect 2438 878 2496 890
rect 2438 602 2450 878
rect 2484 602 2496 878
rect 2438 590 2496 602
rect 2171 574 2233 586
rect 1552 546 1614 558
<< ndiffc >>
rect 1376 234 1410 360
rect 1472 234 1506 360
rect 1568 234 1602 360
rect 1902 198 1936 324
rect 1998 198 2032 324
rect 2094 198 2128 324
rect 2360 286 2394 412
rect 2448 286 2482 412
<< pdiffc >>
rect 1376 558 1410 834
rect 1472 558 1506 834
rect 1568 558 1602 834
rect 1803 586 1837 862
rect 1899 586 1933 862
rect 1995 586 2029 862
rect 2091 586 2125 862
rect 2187 586 2221 862
rect 2362 602 2396 878
rect 2450 602 2484 878
<< psubdiff >>
rect 1365 18 1389 52
rect 1589 18 1613 52
rect 1889 26 1913 60
rect 2113 26 2137 60
rect 2301 24 2325 58
rect 2525 24 2549 58
<< nsubdiff >>
rect 1888 1042 2136 1043
rect 1364 1034 1612 1035
rect 1364 1000 1413 1034
rect 1560 1000 1612 1034
rect 1888 1008 1937 1042
rect 2084 1008 2136 1042
rect 1888 1007 2136 1008
rect 2300 1040 2548 1041
rect 2300 1006 2349 1040
rect 2496 1006 2548 1040
rect 2300 1005 2548 1006
rect 1364 999 1612 1000
<< psubdiffcont >>
rect 1389 18 1589 52
rect 1913 26 2113 60
rect 2325 24 2525 58
<< nsubdiffcont >>
rect 1413 1000 1560 1034
rect 1937 1008 2084 1042
rect 2349 1006 2496 1040
<< poly >>
rect 1320 942 1520 958
rect -288 556 -230 932
rect 1320 908 1338 942
rect 1372 920 1520 942
rect 1852 948 2168 976
rect 1852 946 2172 948
rect 1372 908 1456 920
rect 1320 890 1456 908
rect 1852 900 1884 946
rect 1416 872 1456 890
rect 1426 846 1456 872
rect 1522 846 1552 876
rect 1853 874 1883 900
rect 1949 874 1979 904
rect 2045 874 2075 900
rect 2136 892 2172 946
rect 2141 874 2171 892
rect 2408 890 2438 916
rect -290 460 -116 556
rect 1853 550 1883 574
rect 1044 450 1174 522
rect 1426 372 1456 546
rect 1522 372 1552 546
rect 1734 510 1802 526
rect 1734 476 1752 510
rect 1786 506 1802 510
rect 1846 506 1888 550
rect 1949 548 1979 574
rect 2045 550 2075 574
rect 2044 548 2076 550
rect 2141 548 2171 574
rect 2408 572 2438 590
rect 1786 476 1888 506
rect 1948 504 2076 548
rect 1734 458 1888 476
rect 1738 448 1888 458
rect 1950 388 1988 504
rect 2140 468 2172 548
rect 2406 530 2438 572
rect 2306 514 2438 530
rect 2306 480 2324 514
rect 2358 480 2438 514
rect 2140 392 2178 468
rect 2306 462 2438 480
rect 2308 458 2438 462
rect 2406 446 2438 458
rect 2406 424 2436 446
rect 1822 360 1988 388
rect 2048 362 2178 392
rect 1822 358 1982 360
rect 1822 348 1862 358
rect 1746 288 1862 348
rect 1952 336 1982 358
rect 2048 336 2078 362
rect 1746 254 1764 288
rect 1798 254 1862 288
rect 1746 234 1862 254
rect 1426 196 1456 222
rect 1522 204 1552 222
rect 1522 166 1560 204
rect 2406 248 2436 274
rect 1500 150 1568 166
rect 1952 160 1982 186
rect 2048 160 2078 186
rect 1500 116 1518 150
rect 1552 116 1568 150
rect 1500 98 1568 116
<< polycont >>
rect 1338 908 1372 942
rect 1752 476 1786 510
rect 2324 480 2358 514
rect 1764 254 1798 288
rect 1518 116 1552 150
<< locali >>
rect 1879 1047 2145 1050
rect 1355 1039 1621 1042
rect 1355 996 1361 1039
rect 1616 996 1621 1039
rect 1879 1004 1885 1047
rect 2140 1004 2145 1047
rect 1879 1000 2145 1004
rect 2291 1045 2557 1048
rect 2291 1002 2297 1045
rect 2552 1002 2557 1045
rect 2291 998 2557 1002
rect 1355 992 1621 996
rect 1326 942 1384 958
rect 1326 908 1338 942
rect 1372 908 1384 942
rect 1326 890 1384 908
rect 2362 878 2396 894
rect 1803 862 1837 878
rect 1376 834 1410 850
rect 1376 542 1410 558
rect 1472 834 1506 850
rect 1472 542 1506 558
rect 1568 834 1602 850
rect 1803 570 1837 586
rect 1899 862 1933 878
rect 1899 570 1933 586
rect 1995 862 2029 878
rect 1995 570 2029 586
rect 2091 862 2125 878
rect 2091 570 2125 586
rect 2187 862 2221 878
rect 2362 586 2396 602
rect 2450 878 2484 894
rect 2450 586 2484 602
rect 2187 570 2221 586
rect 1568 542 1602 558
rect 1740 510 1798 526
rect 1740 476 1752 510
rect 1786 476 1798 510
rect 1740 458 1798 476
rect 2312 514 2370 530
rect 2312 480 2324 514
rect 2358 480 2370 514
rect 2312 462 2370 480
rect 2360 412 2394 428
rect 1376 360 1410 376
rect 1376 218 1410 234
rect 1472 360 1506 376
rect 1472 218 1506 234
rect 1568 360 1602 376
rect 1902 324 1936 340
rect 1752 288 1810 304
rect 1752 254 1764 288
rect 1798 254 1810 288
rect 1752 236 1810 254
rect 1568 218 1602 234
rect 1902 182 1936 198
rect 1998 324 2032 340
rect 1998 182 2032 198
rect 2094 324 2128 340
rect 2360 270 2394 286
rect 2448 412 2482 428
rect 2448 270 2482 286
rect 2094 182 2128 198
rect 1506 150 1564 166
rect 1506 116 1518 150
rect 1552 116 1564 150
rect 1506 98 1564 116
<< viali >>
rect 1361 1034 1616 1039
rect 1361 1000 1413 1034
rect 1413 1000 1560 1034
rect 1560 1000 1616 1034
rect 1361 996 1616 1000
rect 1885 1042 2140 1047
rect 1885 1008 1937 1042
rect 1937 1008 2084 1042
rect 2084 1008 2140 1042
rect 1885 1004 2140 1008
rect 2297 1040 2552 1045
rect 2297 1006 2349 1040
rect 2349 1006 2496 1040
rect 2496 1006 2552 1040
rect 2297 1002 2552 1006
rect 1338 908 1372 942
rect 1376 558 1410 834
rect 1472 558 1506 834
rect 1568 558 1602 834
rect 1803 586 1837 862
rect 1899 586 1933 862
rect 1995 586 2029 862
rect 2091 586 2125 862
rect 2187 586 2221 862
rect 2362 602 2396 878
rect 2450 602 2484 878
rect 1752 476 1786 510
rect 2324 480 2358 514
rect 1376 234 1410 360
rect 1472 234 1506 360
rect 1568 234 1602 360
rect 1764 254 1798 288
rect 1902 198 1936 324
rect 1998 198 2032 324
rect 2094 198 2128 324
rect 2360 286 2394 412
rect 2448 286 2482 412
rect 1518 116 1552 150
rect 1886 60 2141 65
rect 1362 52 1617 57
rect 1362 18 1389 52
rect 1389 18 1589 52
rect 1589 18 1617 52
rect 1886 26 1913 60
rect 1913 26 2113 60
rect 2113 26 2141 60
rect 1886 22 2141 26
rect 2298 58 2553 63
rect 2298 24 2325 58
rect 2325 24 2525 58
rect 2525 24 2553 58
rect 2298 20 2553 24
rect 1362 14 1617 18
<< metal1 >>
rect -272 1051 2554 1064
rect -272 1047 2564 1051
rect -272 1039 1885 1047
rect -272 1010 1361 1039
rect 1349 996 1361 1010
rect 1616 1010 1885 1039
rect 1616 996 1628 1010
rect 1780 1004 1885 1010
rect 2140 1045 2564 1047
rect 2140 1010 2297 1045
rect 2140 1004 2226 1010
rect 1780 1000 2226 1004
rect 1780 998 2152 1000
rect 1780 996 1898 998
rect 1349 990 1628 996
rect -300 952 -234 958
rect -300 900 -294 952
rect -242 900 -234 952
rect -300 892 -234 900
rect 1318 952 1388 958
rect 1318 900 1328 952
rect 1380 900 1388 952
rect 1788 908 1840 996
rect 1892 926 2132 966
rect 1318 892 1388 900
rect 1326 890 1384 892
rect 1786 862 1844 908
rect 1892 872 1940 926
rect 2084 874 2132 926
rect 2182 874 2226 1000
rect 2285 1002 2297 1010
rect 2552 1002 2564 1045
rect 2285 996 2564 1002
rect 2350 878 2402 996
rect 1370 842 1416 846
rect 1346 836 1416 842
rect 1214 828 1280 834
rect 1214 776 1220 828
rect 1272 776 1280 828
rect 1346 784 1356 836
rect 1408 834 1416 836
rect 1346 776 1376 784
rect 1214 768 1280 776
rect 1370 628 1376 776
rect 1268 618 1336 624
rect 1268 566 1278 618
rect 1330 566 1336 618
rect 1268 558 1336 566
rect 468 510 542 518
rect 468 458 474 510
rect 526 458 542 510
rect 468 446 542 458
rect 924 508 1106 524
rect 924 456 976 508
rect 1028 456 1106 508
rect 924 450 1106 456
rect 1272 512 1336 558
rect 1364 558 1376 628
rect 1410 558 1416 834
rect 1364 546 1416 558
rect 1466 834 1512 846
rect 1466 558 1472 834
rect 1506 558 1512 834
rect 1364 540 1414 546
rect 930 444 1100 450
rect 930 442 1012 444
rect 1272 378 1344 512
rect 1466 504 1512 558
rect 1562 834 1608 846
rect 1562 558 1568 834
rect 1602 622 1608 834
rect 1640 834 1712 840
rect 1786 838 1803 862
rect 1640 782 1650 834
rect 1702 782 1712 834
rect 1640 774 1712 782
rect 1602 616 1636 622
rect 1628 564 1636 616
rect 1602 558 1636 564
rect 1562 556 1636 558
rect 1664 620 1712 774
rect 1562 546 1608 556
rect 1466 484 1574 504
rect 1466 428 1486 484
rect 1548 428 1574 484
rect 1466 414 1574 428
rect 1272 372 1414 378
rect 1272 360 1416 372
rect 484 290 550 296
rect -100 168 -48 276
rect 484 238 490 290
rect 542 238 550 290
rect 484 230 550 238
rect 1272 234 1376 360
rect 1410 234 1416 360
rect 1272 222 1416 234
rect 1466 360 1512 414
rect 1562 370 1608 372
rect 1664 370 1704 620
rect 1797 586 1803 838
rect 1837 838 1844 862
rect 1893 862 1939 872
rect 1837 586 1843 838
rect 1797 574 1843 586
rect 1893 586 1899 862
rect 1933 586 1939 862
rect 1893 574 1939 586
rect 1989 862 2035 874
rect 1989 586 1995 862
rect 2029 586 2035 862
rect 1989 584 2035 586
rect 2085 862 2131 874
rect 2085 586 2091 862
rect 2125 586 2131 862
rect 1988 532 2038 584
rect 2085 574 2131 586
rect 2181 862 2227 874
rect 2181 586 2187 862
rect 2221 586 2227 862
rect 2350 676 2362 878
rect 2356 602 2362 676
rect 2396 602 2402 878
rect 2356 590 2402 602
rect 2444 878 2490 890
rect 2444 602 2450 878
rect 2484 842 2490 878
rect 2484 836 2544 842
rect 2536 784 2544 836
rect 2484 776 2544 784
rect 2484 736 2490 776
rect 2484 602 2502 736
rect 2444 590 2502 602
rect 2181 574 2227 586
rect 1732 518 1806 526
rect 1732 466 1738 518
rect 1790 466 1806 518
rect 1988 500 2042 532
rect 2188 516 2370 532
rect 2188 500 2240 516
rect 1732 454 1806 466
rect 1986 464 2240 500
rect 2292 514 2370 516
rect 2292 480 2324 514
rect 2358 480 2370 514
rect 2292 464 2370 480
rect 1986 458 2370 464
rect 1986 452 2364 458
rect 1986 450 2276 452
rect 1986 446 2274 450
rect 1466 234 1472 360
rect 1506 234 1512 360
rect 1466 222 1512 234
rect 1560 360 1704 370
rect 1560 234 1568 360
rect 1602 234 1704 360
rect 1988 426 2042 446
rect 1896 324 1942 336
rect 1750 300 1816 306
rect 1750 248 1756 300
rect 1808 248 1816 300
rect 1750 240 1816 248
rect 1752 236 1810 240
rect 1560 222 1704 234
rect 1664 216 1704 222
rect 1896 202 1902 324
rect 1878 198 1902 202
rect 1936 198 1942 324
rect 1988 324 2038 426
rect 2450 424 2502 590
rect 2350 412 2402 424
rect 1988 316 1998 324
rect 1878 186 1942 198
rect 1992 198 1998 316
rect 2032 198 2038 324
rect 1992 186 2038 198
rect 2088 324 2134 336
rect 2088 198 2094 324
rect 2128 198 2134 324
rect 2088 194 2134 198
rect 2350 286 2360 412
rect 2394 286 2402 412
rect -100 120 202 168
rect -96 92 202 120
rect 1500 160 1570 166
rect 1500 108 1510 160
rect 1562 108 1570 160
rect 1500 100 1570 108
rect 1506 98 1564 100
rect 1878 71 1936 186
rect 2086 71 2152 194
rect 728 60 872 62
rect 728 58 886 60
rect 1348 58 1640 68
rect 1874 65 2153 71
rect 2350 69 2402 286
rect 2442 412 2502 424
rect 2442 286 2448 412
rect 2482 356 2502 412
rect 2482 286 2488 356
rect 2442 274 2488 286
rect 1812 58 1886 65
rect -264 57 1886 58
rect -264 14 1362 57
rect 1617 22 1886 57
rect 2141 58 2195 65
rect 2286 63 2565 69
rect 2286 58 2298 63
rect 2141 22 2298 58
rect 1617 20 2298 22
rect 2553 20 2565 63
rect 1617 14 2565 20
rect -264 10 2558 14
rect 1350 8 1629 10
rect 1812 6 1997 10
rect 2028 6 2195 10
<< via1 >>
rect -294 900 -242 952
rect 1328 942 1380 952
rect 1328 908 1338 942
rect 1338 908 1372 942
rect 1372 908 1380 942
rect 1328 900 1380 908
rect 1220 776 1272 828
rect 1356 834 1408 836
rect 1356 784 1376 834
rect 1376 784 1408 834
rect 1278 566 1330 618
rect 474 458 526 510
rect 976 456 1028 508
rect 1650 782 1702 834
rect 1576 564 1602 616
rect 1602 564 1628 616
rect 1486 428 1548 484
rect 490 238 542 290
rect 2484 784 2536 836
rect 1738 510 1790 518
rect 1738 476 1752 510
rect 1752 476 1786 510
rect 1786 476 1790 510
rect 1738 466 1790 476
rect 2240 464 2292 516
rect 1756 288 1808 300
rect 1756 254 1764 288
rect 1764 254 1798 288
rect 1798 254 1808 288
rect 1756 248 1808 254
rect 1510 150 1562 160
rect 1510 116 1518 150
rect 1518 116 1552 150
rect 1552 116 1562 150
rect 1510 108 1562 116
<< metal2 >>
rect 22 964 1738 968
rect -310 962 1738 964
rect -310 952 2624 962
rect -310 900 -294 952
rect -242 900 1328 952
rect 1380 900 2624 952
rect -310 884 2624 900
rect 22 882 2624 884
rect 1298 880 2624 882
rect 1298 878 1732 880
rect 1642 846 2550 850
rect 378 828 1286 842
rect 378 776 1220 828
rect 1272 776 1286 828
rect 378 762 1286 776
rect 1336 836 2550 846
rect 1336 784 1356 836
rect 1408 834 2484 836
rect 1408 784 1650 834
rect 1336 782 1650 784
rect 1702 784 2484 834
rect 2536 784 2550 836
rect 1702 782 2550 784
rect 1336 774 2550 782
rect 1642 770 2550 774
rect -322 540 72 628
rect 1264 618 1638 628
rect 1264 566 1278 618
rect 1330 616 1638 618
rect 1330 566 1576 616
rect 1264 564 1576 566
rect 1628 564 1638 616
rect 1264 550 1638 564
rect 1264 530 1336 550
rect 410 510 538 518
rect 410 458 474 510
rect 526 458 538 510
rect 410 396 538 458
rect 956 508 1336 530
rect 956 456 976 508
rect 1028 456 1336 508
rect 1674 518 1802 526
rect 1674 496 1738 518
rect 956 438 1336 456
rect 1264 436 1336 438
rect 1468 484 1738 496
rect 1468 428 1486 484
rect 1548 466 1738 484
rect 1790 466 1802 518
rect 1548 428 1802 466
rect 2220 516 2596 538
rect 2220 464 2240 516
rect 2292 464 2596 516
rect 2220 446 2596 464
rect 1468 416 1802 428
rect 1674 404 1802 416
rect -304 300 2616 310
rect -304 290 1756 300
rect -304 238 490 290
rect 542 248 1756 290
rect 1808 248 2616 300
rect 542 238 2616 248
rect -304 220 2616 238
rect 1490 166 1578 170
rect 1278 160 1710 166
rect 1278 150 1510 160
rect 22 108 1510 150
rect 1562 108 1710 160
rect 22 90 1710 108
rect 1278 86 1710 90
use dpg2  dpg2_0
timestamp 1710356038
transform 1 0 64 0 1 -46
box -64 46 404 1109
use inv  inv_0
timestamp 1710275825
transform 1 0 1000 0 1 6
box 0 0 320 1063
use inv  inv_1
timestamp 1710275825
transform 1 0 -278 0 1 8
box 0 0 320 1063
use nor  nor_0 nor
timestamp 1710356038
transform 1 0 924 0 1 -58
box -646 56 86 1129
use via_m1_p#0  via_m1_p_0
timestamp 1646951168
transform 1 0 1042 0 1 454
box 0 0 68 68
use via_m1_p#0  via_m1_p_1
timestamp 1646951168
transform 1 0 -304 0 1 886
box 0 0 68 68
<< labels >>
rlabel nwell 621 996 876 1039 1 V
rlabel metal2 2292 446 2596 538 1 Q
rlabel metal1 125 10 325 44 1 GND
rlabel metal2 -322 540 72 628 1 D
rlabel poly -288 460 -230 932 1 clk
rlabel metal2 -304 220 490 310 1 R
rlabel space 14 90 1510 150 1 nclk
<< end >>
