magic
tech sky130A
magscale 1 2
timestamp 1710263695
<< nwell >>
rect -160 170 160 188
rect -161 160 160 170
rect -161 -22 161 160
rect -162 -178 161 -22
rect -162 -190 160 -178
<< pmos >>
rect -63 -150 -33 150
rect 33 -150 63 150
<< pdiff >>
rect -125 138 -63 150
rect -125 -138 -113 138
rect -79 -138 -63 138
rect -125 -150 -63 -138
rect -33 138 33 150
rect -33 -138 -17 138
rect 17 -138 33 138
rect -33 -150 33 -138
rect 63 138 125 150
rect 63 -138 79 138
rect 113 -138 125 138
rect 63 -150 125 -138
<< pdiffc >>
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
<< poly >>
rect -63 150 -33 176
rect 33 150 63 180
rect -63 -178 -33 -150
rect 33 -176 63 -150
<< locali >>
rect -113 138 -79 154
rect -113 -154 -79 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 79 138 113 154
rect 79 -154 113 -138
<< viali >>
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
<< metal1 >>
rect -119 138 -73 150
rect -119 -138 -113 138
rect -79 -138 -73 138
rect -119 -150 -73 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 73 138 119 150
rect 73 -138 79 138
rect 113 -138 119 138
rect 73 -150 119 -138
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
