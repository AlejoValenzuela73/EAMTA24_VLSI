magic
tech sky130A
magscale 1 2
timestamp 1709763159
<< nmos >>
rect -63 -75 -33 75
rect 33 -75 63 75
<< ndiff >>
rect -125 63 -63 75
rect -125 -63 -113 63
rect -79 -63 -63 63
rect -125 -75 -63 -63
rect -33 63 33 75
rect -33 -63 -17 63
rect 17 -63 33 63
rect -33 -75 33 -63
rect 63 63 125 75
rect 63 -63 79 63
rect 113 -63 125 63
rect 63 -75 125 -63
<< ndiffc >>
rect -113 -63 -79 63
rect -17 -63 17 63
rect 79 -63 113 63
<< poly >>
rect -248 152 -34 182
rect -246 145 -34 152
rect -246 111 -215 145
rect -181 124 -34 145
rect -181 116 -33 124
rect -181 111 -152 116
rect -246 90 -152 111
rect -82 100 -33 116
rect -63 75 -33 100
rect 32 92 66 124
rect 33 75 63 92
rect -246 -95 -156 -76
rect -246 -129 -221 -95
rect -187 -129 -156 -95
rect -63 -102 -33 -75
rect 33 -97 63 -75
rect -246 -147 -156 -129
rect -247 -152 -156 -147
rect 32 -152 63 -97
rect -247 -158 63 -152
rect -248 -188 63 -158
<< polycont >>
rect -215 111 -181 145
rect -221 -129 -187 -95
<< locali >>
rect -231 111 -215 145
rect -181 111 -165 145
rect -113 63 -79 79
rect -113 -79 -79 -63
rect -17 63 17 79
rect -17 -79 17 -63
rect 79 63 113 79
rect 79 -79 113 -63
rect -237 -129 -221 -95
rect -187 -129 -171 -95
<< viali >>
rect -215 111 -181 145
rect -113 -63 -79 63
rect -17 -63 17 63
rect 79 -63 113 63
rect -221 -129 -187 -95
<< metal1 >>
rect -298 145 -164 166
rect -298 111 -215 145
rect -181 111 -164 145
rect -298 98 -164 111
rect -119 63 -73 75
rect -119 -63 -113 63
rect -79 -63 -73 63
rect -119 -75 -73 -63
rect -23 63 23 75
rect -23 -63 -17 63
rect 17 -63 23 63
rect -23 -75 23 -63
rect 73 63 119 75
rect 73 -63 79 63
rect 113 -63 119 63
rect 73 -75 119 -63
rect -233 -90 -175 -89
rect -290 -95 -168 -90
rect -290 -129 -221 -95
rect -187 -129 -168 -95
rect -290 -144 -168 -129
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.75 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
